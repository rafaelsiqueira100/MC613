library ieee;
use ieee.std_logic_1164.all;

entity d5to32 is
	port(
		data_in: std_logic_vector (4 downto 0);
		enable: in std_logic;
		data_out: out std_logic_vector (31 downto 0)
	);
end entity;
	
architecture arc of d5to32 is
		signal auxiliar: std_logic_vector(5 downto 0);
begin
	auxiliar <= data_in & enable;
	with auxiliar select
		data_out <= "00000000000000000000000000000001" when "000001",
						"00000000000000000000000000000010" when "100001",
						"00000000000000000000000000000100" when "010001",
						"00000000000000000000000000001000" when "110001",
						"00000000000000000000000000010000" when "001001",
						"00000000000000000000000000100000" when "101001",
						"00000000000000000000000001000000" when "011001",
						"00000000000000000000000010000000" when "111001",
						"00000000000000000000000100000000" when "000101",
						"00000000000000000000001000000000" when "100101",
						"00000000000000000000010000000000" when "010101",
						"00000000000000000000100000000000" when "110101",
						"00000000000000000001000000000000" when "001101",
						"00000000000000000010000000000000" when "101101",
						"00000000000000000100000000000000" when "011101",
						"00000000000000001000000000000000" when "111101",
						"00000000000000010000000000000000" when "000011",
						"00000000000000100000000000000000" when "100011",
						"00000000000001000000000000000000" when "010011",
						"00000000000010000000000000000000" when "110011",
						"00000000000100000000000000000000" when "001011",
						"00000000001000000000000000000000" when "101011",
						"00000000010000000000000000000000" when "011011",
						"00000000100000000000000000000000" when "111011",
						"00000001000000000000000000000000" when "000011",
						"00000010000000000000000000000000" when "100011",
						"00000100000000000000000000000000" when "010011",
						"00001000000000000000000000000000" when "110011",
						"00010000000000000000000000000000" when "001011",
						"00100000000000000000000000000000" when "101011",
						"01000000000000000000000000000000" when "011011",
						"10000000000000000000000000000000" when "111011",
						"00000000000000000000000000000000" when others;
end arc;