<!DOCTYPE html>
<html dir="ltr" class="W0dUmf zIKt9b" lang="pt-BR"><head>
<meta http-equiv="content-type" content="text/html; charset=UTF-8"><!-- base href="https://classroom.google.com/" --><meta name="referrer" content="origin"><meta name="viewport" content="width=device-width, initial-scale=1"><meta name="mobile-web-app-capable" content="yes"><meta name="apple-mobile-web-app-capable" content="yes"><meta name="application-name" content="Google Classroom"><meta name="apple-mobile-web-app-title" content="Google Classroom"><meta name="apple-mobile-web-app-status-bar-style" content="black"><meta name="msapplication-tap-highlight" content="no"><link rel="manifest" crossorigin="use-credentials" href="https://classroom.google.com/_/ClassroomUi/manifest.json"><link rel="home" href="https://classroom.google.com/?lfhs=2"><link rel="msapplication-starturl" href="https://classroom.google.com/?lfhs=2"><link rel="apple-touch-icon-precomposed" href="https://ssl.gstatic.com/classroom/ic_product_classroom_32.png" sizes="32x32"><link rel="msapplication-square32x32logo" href="https://ssl.gstatic.com/classroom/ic_product_classroom_32.png" sizes="32x32"><link rel="apple-touch-icon-precomposed" href="https://ssl.gstatic.com/classroom/ic_product_classroom_48.png" sizes="48x48"><link rel="msapplication-square48x48logo" href="https://ssl.gstatic.com/classroom/ic_product_classroom_48.png" sizes="48x48"><link rel="apple-touch-icon-precomposed" href="https://ssl.gstatic.com/classroom/ic_product_classroom_96.png" sizes="96x96"><link rel="msapplication-square96x96logo" href="https://ssl.gstatic.com/classroom/ic_product_classroom_96.png" sizes="96x96"><link rel="apple-touch-icon-precomposed" href="https://ssl.gstatic.com/classroom/ic_product_classroom_144.png" sizes="144x144"><link rel="msapplication-square144x144logo" href="https://ssl.gstatic.com/classroom/ic_product_classroom_144.png" sizes="144x144"><script src="dec2_to_4_files/cb=gapi.loaded_1" nonce="" async=""></script><script src="dec2_to_4_files/cb=gapi.loaded_0" nonce="" async=""></script><script data-id="_gd" nonce="">window.WIZ_global_data = {"DpimGf":false,"EP1ykd":["/_/*"],"FdrFJe":"-7660840398983927425","Im6cmf":"/_/ClassroomUi","LVIXXb":1,"LoQv7e":false,"MT7f9b":[],"MuJWjd":false,"Pttpvd":"https://connect.corp.google.com/","QrtxK":"0","S06Grb":"112038394563442416565","SNlM0e":"AD_W2oNDbjunZECTRIvwJkg1TSsp:1679956297868","W3Yyqf":"112038394563442416565","WZsZ1e":"M0vAhOfGDwthpy_7/AbZEX3tsZXsLiYaUJ","Yllh3e":"%.@.1679956297702249,180638663,772779554]","YlwcZe":"%.@.3,[1],[3600],2,[15,4,13,14,12,2]]","cfb2h":"boq_apps-edu-classroom-ui_20230313.07_p2","eQxUid":false,"eptZe":"/_/ClassroomUi/","fPDxwd":[1763433,1772879,45814370,47893265,47977019,48410021,48504704,48577232,48642514],"fX0NEc":"%.@.]","gGcLoe":false,"khbx6e":false,"nQyAE":{"Cq67kd":"false","wKmy3":"false","LUVRSd":"false","KfdDpc":"false","wvFeYd":"https://people-pa.googleapis.com/$discovery/rest?version\u003dv2","Ys7BHf":"false","duuZ1c":"true","piHgrf":"false","arUahf":"false","Xr9Q1e":"true","yKLihb":"false","WJMzId":"false","G892ad":"false","xmeGFd":"true","dYFpCd":"false","GFLFFc":"false","ifCQkd":"false","HboSu":"false","sDonxd":"false","L1Y4vd":"false","oC4WDe":"true","votR5b":"false","UvZcsc":"true","qivG0c":"true","eDFRAc":"false","w4j9w":"false","ZyMsw":"false","DTwAnd":"false","JYPDgf":"false","d6y8ud":"false","S60lQe":"false","eyYkRb":"false","ZREghd":"false","WvnWb":"false","X1UVLd":"false","NwDvqe":"false","lW9rfc":"false","RKg7re":"true","D1bn1b":"false"},"oPEP7c":"r243360@dac.unicamp.br","qDCSke":"112038394563442416565","qwAQke":"ClassroomUi","rtQCxc":180,"u9xrGb":"%.@.\"https://drive.google.com/picker\",null,null,null,null,null,null,null,null,null,null,null,[null,null,\"CIvF_fKU_f0CFcdTxAodIq4PLg\",1679956297867986,[48475730,48532127,48545168,48548282,45826083,47809549,48642514,47930869,47809351,1787118,47977019,48494755,47893265,47988271,1714246,45814370,47856925,47835375,47860858,1772879,47948077,45754602,45686039,48638933,45775441,1773158,1706538,1729889,48577232,48504704,47807826,48539282,48511759,45771378,1763433,45758671,45774183,48663492,47790498,45735197,48573003,47844885,48410021,49617885,49365716,48475720,48532116,48545154,48548272,45826071,47930858,47809341,48494744,47893254,47988260,47856911,47835361,47948067,45754588,48638923,47807816,48511749,45774169,48663482,47790484,48572993,47844875,49617874,49365706],2],null,null,1000,\"\",null,null,[null,null,\"p\",1800000,null,null,null,10000,39000,120000,2,null,100,3100,null,\"/punctual/prod/homeroom_prod\"],null,null,null,null,null,null,[null,null,\"https://gstatic.com/classroom/themes/img_backtoschool.jpg\"],null,\"r\",null,null,null,\"\",0,null,null,null,null,null,null,null,10,null,null,5,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,10,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,true,null,null,null,null,null,null,null,null,null,null,20,null,null,null,null,null,null,null,null,1000,null,null,\"{size}\",20,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,\"https://calendar.google.com\",null,null,null,[100,604800000,2,0.5],null,null,null,null,null,null,null,null,null,null,null,null,null,20,null,null,null,\"AIzaSyAewGK8j9KoyT94rEj-weBpysMvzMQzGvk\",\"https://www.googleapis.com/drive/v2internal\",null,null,null,null,null,false,null,null,null,true,true,null,null,null,null,null,null,null,null,null,null,null,null,\"https://docs.google.com\",\"https://drive.google.com\",null,100,null,null,null,null,true,null,\"unicamp.br\",\"^video/|^application/(x-flash-video|vnd\\\\.google-apps\\\\.video|video)$|^application/vnd\\\\.google-apps\\\\.drive-sdk\\\\.\",null,null,null,null,\"https://lh3.googleusercontent.com/a/default-user\\u003ds72-c-fbw\\u003d1\",null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,15,null,null,false,null,null,null,null,null,null,false,null,null,null,null,null,null,null,null,null,null,null,null,null,300000,null,null,null,null,null,null,null,10,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,\"//ssl.gstatic.com/classroom/favicon.png\",null,\"30751363934\",\"https://classroom.google.com/\",null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,true,null,null,null,4000,1.3,null,null,false,null,[3],null,null,null,null,null,null,null,null,null,null,null,true,null,null,null,null,true,false,null,null,null,null,null,true,null,null,null,null,null,[true,\"96485\",\"AIzaSyBqt2sx2fvfwP502G4u_Mu_kRmei_3A2OU\",null,false],null,null,null,null,null,false,null,false,null,null,null,null,null,null,null,null,null,200,null,null,null,null,null,null,null,null,null,false,null,null,null,null,null,null,false,null,null,null,null,true,null,null,true,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,true,\"BR\",null,null,null,null,null,null,[\"https://workspace.google.com\"],null,null,null,null,[false,null,null,null,null,null,null,false,false],null,null,null,null,null,false,null,null,1,null,null,null,false,null,null,null,null,null,null,null,null,null,null,false,null,false,null,1800000,null,null,false,null,null,null,[false,null,[null,null,null,\"https://classroom.google.com/ps/create\"],true,true],730,null,false,false,false,true,true,false,true,false,false,false,false,false,false,false,false,false,false,false,false]","vLjptb":"112038394563442416565","w2btAe":"%.@.\"112038394563442416565\",\"112038394563442416565\",\"0\",false,null,null,true,false]","x3UoP":"%.@.[\"30751363934\"],\"Rafael Andre Alves De Siqueira\",\"r243360@dac.unicamp.br\",[null,[6,12,48,46,56,61,67,73,87,83],null,1,3,2,null,null,true,false],\"//lh3.googleusercontent.com/a/AGNmyxbGKcB41E-oqOD3N45dzBlNoIb7BH01Q9jZOZNGSA\",3,1637183191240,null,false,\"Rafael Andre Alves De Siqueira r243360@dac.unicamp.br\",1,\"Rafael Andre Alves De Siqueira r243360@dac.unicamp.br\",\"Andre Alves De Siqueira Rafael r243360@dac.unicamp.br\",false,false,1,null,null,null,null,[1,\"unicamp.br\",2],true,null,null,null,true,true,false]","x7Mded":"%.@.1,null,300,75,true]","zChJod":"%.@.]"};</script><script nonce="">(function(){'use strict';var a=window,d=a.performance,l=k();a.cc_latency_start_time=d&&d.now?0:d&&d.timing&&d.timing.navigationStart?d.timing.navigationStart:l;function k(){return d&&d.now?d.now():(new Date).getTime()}function n(e){if(d&&d.now&&d.mark){var g=d.mark(e);if(g)return g.startTime;if(d.getEntriesByName&&(e=d.getEntriesByName(e).pop()))return e.startTime}return k()}a.onaft=function(){n("aft")};a._isLazyImage=function(e){return e.hasAttribute("data-src")||e.hasAttribute("data-ils")||"lazy"===e.getAttribute("loading")};
a.l=function(e){function g(b){var c={};c[b]=k();a.cc_latency.push(c)}function m(b){var c=n("iml");b.setAttribute("data-iml",c);return c}a.cc_aid=e;a.iml_start=a.cc_latency_start_time;a.css_size=0;a.cc_latency=[];a.ccTick=g;a.onJsLoad=function(){g("jsl")};a.onCssLoad=function(){g("cssl")};a._isVisible=function(b,c){if(!c||"none"==c.style.display)return!1;var f=b.defaultView;if(f&&f.getComputedStyle&&(f=f.getComputedStyle(c),"0px"==f.height||"0px"==f.width||"hidden"==f.visibility))return!1;if(!c.getBoundingClientRect)return!0;
var h=c.getBoundingClientRect();c=h.left+a.pageXOffset;f=h.top+a.pageYOffset;if(0>f+h.height||0>c+h.width||0>=h.height||0>=h.width)return!1;b=b.documentElement;return f<=(a.innerHeight||b.clientHeight)&&c<=(a.innerWidth||b.clientWidth)};a._recordImlEl=m;document.documentElement.addEventListener("load",function(b){b=b.target;var c;"IMG"!=b.tagName||b.hasAttribute("data-iid")||a._isLazyImage(b)||b.hasAttribute("data-noaft")||(c=m(b));if(a.aft_counter&&(b=a.aft_counter.indexOf(b),-1!==b&&(b=1===a.aft_counter.splice(b,
1).length,0===a.aft_counter.length&&b&&c)))a.onaft(c)},!0);a.prt=-1;a.wiz_tick=function(){var b=n("prt");a.prt=b}};}).call(this);
l('qenh')</script><script nonce="">var _F_cssRowKey = 'boq-apps-edu.ClassroomUi.TtUpWVPKfDY.L.F4.O';var _F_combinedSignature = 'AGEDDAu0O65YApLIV9RqhianbMeIWHpdUg';function _DumpException(e) {throw e;}</script><style data-href="https://www.gstatic.com/_/mss/boq-apps-edu/_/ss/k=boq-apps-edu.ClassroomUi.TtUpWVPKfDY.L.F4.O/am=BHgWAgAC/d=1/ed=1/rs=AGEDDAsCoucIn376zTYuTYouSXkzYy6Fyg/m=streamview,_b,_tp,_r" nonce="">@keyframes mdc-ripple-fg-radius-in{0%{animation-timing-function:cubic-bezier(0.4,0,0.2,1);transform:translate(var(--mdc-ripple-fg-translate-start,0)) scale(1)}to{transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}}@keyframes mdc-ripple-fg-opacity-in{0%{animation-timing-function:linear;opacity:0}to{opacity:var(--mdc-ripple-fg-opacity,0)}}@keyframes mdc-ripple-fg-opacity-out{0%{animation-timing-function:linear;opacity:var(--mdc-ripple-fg-opacity,0)}to{opacity:0}}.VfPpkd-ksKsZd-XxIAqe{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;will-change:transform,opacity;position:relative;outline:none;overflow:hidden}.VfPpkd-ksKsZd-XxIAqe::before,.VfPpkd-ksKsZd-XxIAqe::after{position:absolute;-moz-border-radius:50%;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-ksKsZd-XxIAqe::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-ksKsZd-XxIAqe::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf::after{animation:mdc-ripple-fg-opacity-out 150ms;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-ksKsZd-XxIAqe::before,.VfPpkd-ksKsZd-XxIAqe::after{top:-moz-calc(50% - 100%);top:calc(50% - 100%);left:-moz-calc(50% - 100%);left:calc(50% - 100%);width:200%;height:200%}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded],.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd{overflow:visible}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded]::before,.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded]::after,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::before,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::after{top:-moz-calc(50% - 50%);top:calc(50% - 50%);left:-moz-calc(50% - 50%);left:calc(50% - 50%);width:100%;height:100%}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::before,.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::after,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::before,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::after{top:var(--mdc-ripple-top,calc(50% - 50%));left:var(--mdc-ripple-left,calc(50% - 50%));width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::after,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-ksKsZd-XxIAqe::before,.VfPpkd-ksKsZd-XxIAqe::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-ksKsZd-XxIAqe:hover::before,.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,0.04)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,0.12)}.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d)::after{transition:opacity 150ms linear}.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d):active::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-Bz112c-LgbsSe{font-size:24px;width:48px;height:48px;padding:12px}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:48px;max-width:48px}.VfPpkd-Bz112c-LgbsSe.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:40px;height:40px;margin-top:4px;margin-bottom:4px;margin-right:4px;margin-left:4px}.VfPpkd-Bz112c-LgbsSe.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:40px;max-width:40px}.VfPpkd-Bz112c-LgbsSe:disabled{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-disabled-on-light,rgba(0,0,0,.38))}.VfPpkd-Bz112c-LgbsSe svg,.VfPpkd-Bz112c-LgbsSe img{width:24px;height:24px}.VfPpkd-Bz112c-LgbsSe{display:inline-block;position:relative;-moz-box-sizing:border-box;box-sizing:border-box;border:none;outline:none;background-color:transparent;fill:currentColor;color:inherit;text-decoration:none;cursor:pointer;-moz-user-select:none;user-select:none;z-index:0;overflow:visible}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:48px;left:50%;width:48px;transform:translate(-50%,-50%)}@media screen and (forced-colors:active){.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-J1Ukfc-LhBDec,.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-J1Ukfc-LhBDec{display:block}}.VfPpkd-Bz112c-LgbsSe:disabled{cursor:default;pointer-events:none}.VfPpkd-Bz112c-LgbsSe[hidden]{display:none}.VfPpkd-Bz112c-LgbsSe-OWXEXe-KVuj8d-Q3DXx{-moz-box-align:center;align-items:center;display:-moz-inline-box;display:inline-flex;-moz-box-pack:center;justify-content:center}.VfPpkd-Bz112c-J1Ukfc-LhBDec{pointer-events:none;border:2px solid transparent;border-radius:6px;-moz-box-sizing:content-box;box-sizing:content-box;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:100%;width:100%;display:none}@media screen and (forced-colors:active){.VfPpkd-Bz112c-J1Ukfc-LhBDec{border-color:CanvasText}}.VfPpkd-Bz112c-J1Ukfc-LhBDec::after{content:"";border:2px solid transparent;border-radius:8px;display:block;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-Bz112c-J1Ukfc-LhBDec::after{border-color:CanvasText}}.VfPpkd-Bz112c-kBDsod{display:inline-block}.VfPpkd-Bz112c-kBDsod.VfPpkd-Bz112c-kBDsod-OWXEXe-IT5dJd,.VfPpkd-Bz112c-LgbsSe-OWXEXe-IT5dJd .VfPpkd-Bz112c-kBDsod{display:none}.VfPpkd-Bz112c-LgbsSe-OWXEXe-IT5dJd .VfPpkd-Bz112c-kBDsod.VfPpkd-Bz112c-kBDsod-OWXEXe-IT5dJd{display:inline-block}.VfPpkd-Bz112c-mRLv6{height:100%;left:0;outline:none;position:absolute;top:0;width:100%}.VfPpkd-Bz112c-LgbsSe{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-Bz112c-Jh9lGc::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-Bz112c-Jh9lGc::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-Bz112c-Jh9lGc::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{top:0;left:0;width:100%;height:100%}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0);width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-Bz112c-LgbsSe:hover .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc{height:100%;left:0;pointer-events:none;position:absolute;top:0;width:100%;z-index:-1}.VfPpkd-dgl2Hf-ppHlrf-sM5MNb{display:inline}.VfPpkd-LgbsSe{position:relative;display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center;-moz-box-pack:center;justify-content:center;-moz-box-sizing:border-box;box-sizing:border-box;min-width:64px;border:none;outline:none;line-height:inherit;-moz-user-select:none;user-select:none;-webkit-appearance:none;overflow:visible;vertical-align:middle;background:transparent}.VfPpkd-LgbsSe .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-LgbsSe::-moz-focus-inner{padding:0;border:0}.VfPpkd-LgbsSe:active{outline:none}.VfPpkd-LgbsSe:hover{cursor:pointer}.VfPpkd-LgbsSe:disabled{cursor:default;pointer-events:none}.VfPpkd-LgbsSe[hidden]{display:none}.VfPpkd-LgbsSe .VfPpkd-kBDsod{margin-left:0;margin-right:8px;display:inline-block;position:relative;vertical-align:top}[dir=rtl] .VfPpkd-LgbsSe .VfPpkd-kBDsod,.VfPpkd-LgbsSe .VfPpkd-kBDsod[dir=rtl]{margin-left:8px;margin-right:0}.VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge{font-size:0;position:absolute;transform:translate(-50%,-50%);top:50%;left:50%;line-height:normal}.VfPpkd-LgbsSe .VfPpkd-vQzf8d{position:relative}.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec{pointer-events:none;border:2px solid transparent;border-radius:6px;-moz-box-sizing:content-box;box-sizing:content-box;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px);display:none}@media screen and (forced-colors:active){.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec{border-color:CanvasText}}.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec::after{content:"";border:2px solid transparent;border-radius:8px;display:block;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec::after{border-color:CanvasText}}@media screen and (forced-colors:active){.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-J1Ukfc-LhBDec,.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-J1Ukfc-LhBDec{display:block}}.VfPpkd-LgbsSe .VfPpkd-RLmnJb{position:absolute;top:50%;height:48px;left:0;right:0;transform:translateY(-50%)}.VfPpkd-vQzf8d+.VfPpkd-kBDsod{margin-left:8px;margin-right:0}[dir=rtl] .VfPpkd-vQzf8d+.VfPpkd-kBDsod,.VfPpkd-vQzf8d+.VfPpkd-kBDsod[dir=rtl]{margin-left:0;margin-right:8px}svg.VfPpkd-kBDsod{fill:currentColor}.VfPpkd-LgbsSe-OWXEXe-dgl2Hf{margin-top:6px;margin-bottom:6px}.VfPpkd-LgbsSe{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;text-decoration:none}.VfPpkd-LgbsSe{padding:0 8px 0 8px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ{transition:box-shadow .28s cubic-bezier(.4,0,.2,1);padding:0 16px 0 16px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 12px 0 16px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 16px 0 12px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb{transition:box-shadow .28s cubic-bezier(.4,0,.2,1);padding:0 16px 0 16px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 12px 0 16px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 16px 0 12px}.VfPpkd-LgbsSe-OWXEXe-INsAgc{border-style:solid;transition:border .28s cubic-bezier(.4,0,.2,1)}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc{border-style:solid;border-color:transparent}.VfPpkd-LgbsSe{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{z-index:0}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-Jh9lGc::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-Jh9lGc::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-Jh9lGc::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{top:-50%;left:-50%;width:200%;height:200%}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-Jh9lGc{position:absolute;-moz-box-sizing:content-box;box-sizing:content-box;overflow:hidden;z-index:0;top:0;left:0;bottom:0;right:0}.VfPpkd-LgbsSe{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px}.VfPpkd-LgbsSe:not(:disabled){color:#6200ee}.VfPpkd-LgbsSe:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{background-color:#6200ee}.VfPpkd-LgbsSe:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-text-button-pressed-state-layer-opacity,0.12)}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(:disabled){background-color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:disabled{background-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(:disabled){color:#fff}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc::after{background-color:#fff}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.08}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-filled-button-pressed-state-layer-opacity,0.24)}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px;box-shadow:0 3px 1px -2px rgba(0,0,0,.2),0 2px 2px 0 rgba(0,0,0,.14),0 1px 5px 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled){background-color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled{background-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled){color:#fff}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc::after{background-color:#fff}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.08}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-protected-button-pressed-state-layer-opacity,0.24)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):focus{box-shadow:0 2px 4px -1px rgba(0,0,0,.2),0 4px 5px 0 rgba(0,0,0,.14),0 1px 10px 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:hover{box-shadow:0 2px 4px -1px rgba(0,0,0,.2),0 4px 5px 0 rgba(0,0,0,.14),0 1px 10px 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled):active{box-shadow:0 5px 5px -3px rgba(0,0,0,.2),0 8px 10px 1px rgba(0,0,0,.14),0 3px 14px 2px rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled{box-shadow:0 0 0 0 rgba(0,0,0,.2),0 0 0 0 rgba(0,0,0,.14),0 0 0 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px;padding:0 15px 0 15px;border-width:1px}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(:disabled){color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-INsAgc:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc::after{background-color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-INsAgc:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(:disabled){border-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc:disabled{border-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 11px 0 15px}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 15px 0 11px}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc{top:-1px;left:-1px;bottom:-1px;right:-1px;border-width:1px}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-RLmnJb{left:-1px;width:calc(100% + 2px)}.nCP5yc{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.nCP5yc .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.nCP5yc:not(:disabled){background-color:rgb(26,115,232);background-color:var(--gm-fillbutton-container-color,rgb(26,115,232))}.nCP5yc:not(:disabled){color:#fff;color:var(--gm-fillbutton-ink-color,#fff)}.nCP5yc:disabled{background-color:rgba(60,64,67,.12);background-color:var(--gm-fillbutton-disabled-container-color,rgba(60,64,67,.12))}.nCP5yc:disabled{color:rgba(60,64,67,.38);color:var(--gm-fillbutton-disabled-ink-color,rgba(60,64,67,.38))}.nCP5yc .VfPpkd-Jh9lGc::before,.nCP5yc .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36);background-color:var(--gm-fillbutton-state-color,rgb(32,33,36))}.nCP5yc:hover .VfPpkd-Jh9lGc::before,.nCP5yc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}.nCP5yc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}.nCP5yc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}.nCP5yc .VfPpkd-BFbNVe-bF1uUb{opacity:0}.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#fff}@media (-ms-high-contrast:active),screen and (forced-colors:active){.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.nCP5yc:hover{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-fillbutton-ambientshadow-color,rgba(60,64,67,.15))}.nCP5yc:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.nCP5yc:active{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(60,64,67,.3)),0 2px 6px 2px var(--gm-fillbutton-ambientshadow-color,rgba(60,64,67,.15))}.nCP5yc:active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Rj2Mlf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.Rj2Mlf .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.Rj2Mlf:not(:disabled){color:rgb(26,115,232);color:var(--gm-hairlinebutton-ink-color,rgb(26,115,232))}.Rj2Mlf:not(:disabled){border-color:rgb(218,220,224);border-color:var(--gm-hairlinebutton-outline-color,rgb(218,220,224))}.Rj2Mlf:not(:disabled):hover{border-color:rgb(218,220,224);border-color:var(--gm-hairlinebutton-outline-color,rgb(218,220,224))}.Rj2Mlf:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Rj2Mlf:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(23,78,166);border-color:var(--gm-hairlinebutton-outline-color--stateful,rgb(23,78,166))}.Rj2Mlf:not(:disabled):active,.Rj2Mlf:not(:disabled):focus:active{border-color:rgb(218,220,224);border-color:var(--gm-hairlinebutton-outline-color,rgb(218,220,224))}.Rj2Mlf:disabled{color:rgba(60,64,67,.38);color:var(--gm-hairlinebutton-disabled-ink-color,rgba(60,64,67,.38))}.Rj2Mlf:disabled{border-color:rgba(60,64,67,.12);border-color:var(--gm-hairlinebutton-disabled-outline-color,rgba(60,64,67,.12))}.Rj2Mlf:hover:not(:disabled),.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.Rj2Mlf:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-hairlinebutton-ink-color--stateful,rgb(23,78,166))}.Rj2Mlf .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.Rj2Mlf .VfPpkd-Jh9lGc::before,.Rj2Mlf .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-hairlinebutton-state-color,rgb(26,115,232))}.Rj2Mlf:hover .VfPpkd-Jh9lGc::before,.Rj2Mlf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.b9hyVd{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);border-width:0;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.b9hyVd:not(:disabled){background-color:#fff;background-color:var(--gm-protectedbutton-container-color,#fff)}.b9hyVd:not(:disabled){color:rgb(26,115,232);color:var(--gm-protectedbutton-ink-color,rgb(26,115,232))}.b9hyVd:disabled{background-color:rgba(60,64,67,.12);background-color:var(--gm-protectedbutton-disabled-container-color,rgba(60,64,67,.12))}.b9hyVd:disabled{color:rgba(60,64,67,.38);color:var(--gm-protectedbutton-disabled-ink-color,rgba(60,64,67,.38))}.b9hyVd:hover:not(:disabled),.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.b9hyVd:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-protectedbutton-ink-color--stateful,rgb(23,78,166))}.b9hyVd .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus{border-width:0;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-BFbNVe-bF1uUb,.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd:hover{border-width:0;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 2px 6px 2px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd:not(:disabled):active{border-width:0;box-shadow:0 1px 3px 0 rgba(60,64,67,.3),0 4px 8px 3px rgba(60,64,67,.15);box-shadow:0 1px 3px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 4px 8px 3px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd .VfPpkd-Jh9lGc::before,.b9hyVd .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-protectedbutton-state-color,rgb(26,115,232))}.b9hyVd:hover .VfPpkd-Jh9lGc::before,.b9hyVd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.b9hyVd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.Kjnxrf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.Kjnxrf .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.Kjnxrf:not(:disabled){background-color:rgb(232,240,254)}.Kjnxrf:not(:disabled){color:rgb(25,103,210)}.Kjnxrf:disabled{background-color:rgba(60,64,67,.12)}.Kjnxrf:disabled{color:rgba(60,64,67,.38)}.Kjnxrf:hover:not(:disabled),.Kjnxrf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.Kjnxrf:active:not(:disabled){color:rgb(23,78,166)}.Kjnxrf .VfPpkd-Jh9lGc::before,.Kjnxrf .VfPpkd-Jh9lGc::after{background-color:rgb(25,103,210);background-color:var(--mdc-ripple-color,rgb(25,103,210))}.Kjnxrf:hover .VfPpkd-Jh9lGc::before,.Kjnxrf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.Kjnxrf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.Kjnxrf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.Kjnxrf .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(25,103,210)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.Kjnxrf:hover{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15)}.Kjnxrf:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Kjnxrf:not(:disabled):active{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15)}.Kjnxrf:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.ksBjEc{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none}.ksBjEc .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.ksBjEc:not(:disabled){background-color:transparent}.ksBjEc:not(:disabled){color:rgb(26,115,232);color:var(--gm-colortextbutton-ink-color,rgb(26,115,232))}.ksBjEc:disabled{color:rgba(60,64,67,.38);color:var(--gm-colortextbutton-disabled-ink-color,rgba(60,64,67,.38))}.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.ksBjEc:hover:not(:disabled),.ksBjEc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.ksBjEc:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-colortextbutton-ink-color--stateful,rgb(23,78,166))}.ksBjEc .VfPpkd-Jh9lGc::before,.ksBjEc .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-colortextbutton-state-color,rgb(26,115,232))}.ksBjEc:hover .VfPpkd-Jh9lGc::before,.ksBjEc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.ksBjEc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.ksBjEc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.LjDxcd{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none}.LjDxcd .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.LjDxcd:not(:disabled){color:rgb(95,99,104);color:var(--gm-neutraltextbutton-ink-color,rgb(95,99,104))}.LjDxcd:disabled{color:rgba(60,64,67,.38);color:var(--gm-neutraltextbutton-disabled-ink-color,rgba(60,64,67,.38))}.LjDxcd:hover:not(:disabled),.LjDxcd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.LjDxcd:active:not(:disabled){color:rgb(32,33,36);color:var(--gm-neutraltextbutton-ink-color--stateful,rgb(32,33,36))}.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(95,99,104)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.LjDxcd .VfPpkd-Jh9lGc::before,.LjDxcd .VfPpkd-Jh9lGc::after{background-color:rgb(95,99,104);background-color:var(--gm-neutraltextbutton-state-color,rgb(95,99,104))}.LjDxcd:hover .VfPpkd-Jh9lGc::before,.LjDxcd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.LjDxcd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.LjDxcd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.DuMIQc{padding:0 24px 0 24px}.P62QJc{padding:0 23px 0 23px;border-width:1px}.P62QJc.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 11px 0 23px}.P62QJc.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 23px 0 11px}.P62QJc .VfPpkd-Jh9lGc{top:-1px;left:-1px;bottom:-1px;right:-1px;border-width:1px}.P62QJc .VfPpkd-RLmnJb{left:-1px;width:calc(100% + 2px)}.yHy1rc{z-index:0}.yHy1rc .VfPpkd-Bz112c-Jh9lGc::before,.yHy1rc .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.yHy1rc:disabled{color:rgba(60,64,67,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(60,64,67,.38))}.fzRBVc{z-index:0}.fzRBVc .VfPpkd-Bz112c-Jh9lGc::before,.fzRBVc .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.fzRBVc:disabled{color:rgba(60,64,67,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(60,64,67,.38))}.WpHeLc{height:100%;left:0;position:absolute;top:0;width:100%;outline:none}[dir=rtl] .HDnnrf .VfPpkd-kBDsod,.HDnnrf .VfPpkd-kBDsod[dir=rtl]{transform:scaleX(-1)}[dir=rtl] .QDwDD,.QDwDD[dir=rtl]{transform:scaleX(-1)}.PDpWxe{will-change:unset}.LQeN7 .VfPpkd-J1Ukfc-LhBDec{pointer-events:none;border:2px solid rgb(24,90,188);border-radius:6px;-moz-box-sizing:content-box;box-sizing:content-box;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.LQeN7 .VfPpkd-J1Ukfc-LhBDec{border-color:CanvasText}}.LQeN7 .VfPpkd-J1Ukfc-LhBDec::after{content:"";border:2px solid rgb(232,240,254);border-radius:8px;display:block;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.LQeN7 .VfPpkd-J1Ukfc-LhBDec::after{border-color:CanvasText}}.LQeN7.gmghec .VfPpkd-J1Ukfc-LhBDec{display:inline-block}@media (-ms-high-contrast:active),(-ms-high-contrast:none){.LQeN7.gmghec .VfPpkd-J1Ukfc-LhBDec{display:none}}.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec{pointer-events:none;border:2px solid rgb(24,90,188);border-radius:6px;-moz-box-sizing:content-box;box-sizing:content-box;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:100%;width:100%}@media screen and (forced-colors:active){.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec{border-color:CanvasText}}.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec::after{content:"";border:2px solid rgb(232,240,254);border-radius:8px;display:block;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec::after{border-color:CanvasText}}.mN1ivc.gmghec .VfPpkd-Bz112c-J1Ukfc-LhBDec{display:inline-block}@media (-ms-high-contrast:active),(-ms-high-contrast:none){.mN1ivc.gmghec .VfPpkd-Bz112c-J1Ukfc-LhBDec{display:none}}.MyRpB .VfPpkd-kBDsod,.MyRpB .VfPpkd-vQzf8d{opacity:0}.VfPpkd-MPu53c{padding:11px;padding:calc((var(--mdc-checkbox-ripple-size, 40px) - 18px)/2);margin:0;margin:calc((var(--mdc-checkbox-touch-target-size, 40px) - 40px)/2)}.VfPpkd-MPu53c .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c .VfPpkd-OYHm6b::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-MPu53c:hover .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after{transition:opacity .15s linear}.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:#018786;background-color:var(--mdc-ripple-color,var(--mdc-theme-secondary,#018786))}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:hover .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after{transition:opacity .15s linear}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:#018786;background-color:var(--mdc-ripple-color,var(--mdc-theme-secondary,#018786))}.VfPpkd-MPu53c .VfPpkd-YQoJzd{top:11px;top:calc((var(--mdc-checkbox-ripple-size, 40px) - 18px)/2);left:11px;left:calc((var(--mdc-checkbox-ripple-size, 40px) - 18px)/2)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe{top:0;top:calc((40px - var(--mdc-checkbox-touch-target-size, 40px))/2);right:0;right:calc((40px - var(--mdc-checkbox-touch-target-size, 40px))/2);left:0;left:calc((40px - var(--mdc-checkbox-touch-target-size, 40px))/2);width:40px;width:var(--mdc-checkbox-touch-target-size,40px);height:40px;height:var(--mdc-checkbox-touch-target-size,40px)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgba(0,0,0,.54);border-color:var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54));background-color:transparent}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#018786;border-color:var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786));background-color:#018786;background-color:var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786))}@keyframes mdc-checkbox-fade-in-background-8A000000FF01878600000000FF018786{0%{border-color:rgba(0,0,0,.54);border-color:var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54));background-color:transparent}50%{border-color:#018786;border-color:var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786));background-color:#018786;background-color:var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786))}}@keyframes mdc-checkbox-fade-out-background-8A000000FF01878600000000FF018786{0%,80%{border-color:#018786;border-color:var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786));background-color:#018786;background-color:var(--mdc-checkbox-checked-color,var(--mdc-theme-secondary,#018786))}100%{border-color:rgba(0,0,0,.54);border-color:var(--mdc-checkbox-unchecked-color,rgba(0,0,0,.54));background-color:transparent}}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-8A000000FF01878600000000FF018786}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-8A000000FF01878600000000FF018786}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgba(0,0,0,.38);border-color:var(--mdc-checkbox-disabled-color,rgba(0,0,0,.38));background-color:transparent}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:checked~.VfPpkd-YQoJzd,.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate~.VfPpkd-YQoJzd,.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true][disabled]~.VfPpkd-YQoJzd{border-color:transparent;background-color:rgba(0,0,0,.38);background-color:var(--mdc-checkbox-disabled-color,rgba(0,0,0,.38))}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:#fff;color:var(--mdc-checkbox-ink-color,#fff)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:#fff;border-color:var(--mdc-checkbox-ink-color,#fff)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:#fff;color:var(--mdc-checkbox-ink-color,#fff)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:#fff;border-color:var(--mdc-checkbox-ink-color,#fff)}@keyframes mdc-checkbox-unchecked-checked-checkmark-path{0%,50%{stroke-dashoffset:29.7833385}50%{animation-timing-function:cubic-bezier(0,0,.2,1)}100%{stroke-dashoffset:0}}@keyframes mdc-checkbox-unchecked-indeterminate-mixedmark{0%,68.2%{transform:scaleX(0)}68.2%{animation-timing-function:cubic-bezier(0,0,0,1)}100%{transform:scaleX(1)}}@keyframes mdc-checkbox-checked-unchecked-checkmark-path{from{animation-timing-function:cubic-bezier(.4,0,1,1);opacity:1;stroke-dashoffset:0}to{opacity:0;stroke-dashoffset:-29.7833385}}@keyframes mdc-checkbox-checked-indeterminate-checkmark{from{animation-timing-function:cubic-bezier(0,0,.2,1);transform:rotate(0deg);opacity:1}to{transform:rotate(45deg);opacity:0}}@keyframes mdc-checkbox-indeterminate-checked-checkmark{from{animation-timing-function:cubic-bezier(.14,0,0,1);transform:rotate(45deg);opacity:0}to{transform:rotate(1turn);opacity:1}}@keyframes mdc-checkbox-checked-indeterminate-mixedmark{from{animation-timing-function:mdc-animation-deceleration-curve-timing-function;transform:rotate(-45deg);opacity:0}to{transform:rotate(0deg);opacity:1}}@keyframes mdc-checkbox-indeterminate-checked-mixedmark{from{animation-timing-function:cubic-bezier(.14,0,0,1);transform:rotate(0deg);opacity:1}to{transform:rotate(315deg);opacity:0}}@keyframes mdc-checkbox-indeterminate-unchecked-mixedmark{0%{animation-timing-function:linear;transform:scaleX(1);opacity:1}32.8%,100%{transform:scaleX(0);opacity:0}}.VfPpkd-MPu53c{display:inline-block;position:relative;-moz-box-flex:0;flex:0 0 18px;-moz-box-sizing:content-box;box-sizing:content-box;width:18px;height:18px;line-height:0;white-space:nowrap;cursor:pointer;vertical-align:bottom}.VfPpkd-MPu53c[hidden]{display:none}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec,.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec{pointer-events:none;border:2px solid transparent;border-radius:6px;-moz-box-sizing:content-box;box-sizing:content-box;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:100%;width:100%}@media screen and (forced-colors:active){.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec,.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec{border-color:CanvasText}}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec::after,.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec::after{content:"";border:2px solid transparent;border-radius:8px;display:block;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-sMek6-LhBDec::after,.VfPpkd-MPu53c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-sMek6-LhBDec::after{border-color:CanvasText}}@media (-ms-high-contrast:none){.VfPpkd-MPu53c .VfPpkd-sMek6-LhBDec{display:none}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-SJnn3d{margin:0 1px}}.VfPpkd-MPu53c-OWXEXe-OWB6Me{cursor:default;pointer-events:none}.VfPpkd-YQoJzd{display:-moz-inline-box;display:inline-flex;position:absolute;-moz-box-align:center;align-items:center;-moz-box-pack:center;justify-content:center;-moz-box-sizing:border-box;box-sizing:border-box;width:18px;height:18px;border:2px solid currentColor;border-radius:2px;background-color:transparent;pointer-events:none;will-change:background-color,border-color;transition:background-color 90ms 0ms cubic-bezier(.4,0,.6,1),border-color 90ms 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-HUofsb{position:absolute;top:0;right:0;bottom:0;left:0;width:100%;opacity:0;transition:opacity .18s 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-HUofsb{opacity:1}.VfPpkd-HUofsb-Jt5cK{transition:stroke-dashoffset .18s 0ms cubic-bezier(.4,0,.6,1);stroke:currentColor;stroke-width:3.12px;stroke-dashoffset:29.7833385;stroke-dasharray:29.7833385}.VfPpkd-SJnn3d{width:100%;height:0;transform:scaleX(0) rotate(0deg);border-width:1px;border-style:solid;opacity:0;transition:opacity 90ms 0ms cubic-bezier(.4,0,.6,1),transform 90ms 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-YQoJzd,.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-YQoJzd,.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-YQoJzd,.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-YQoJzd{animation-duration:.18s;animation-timing-function:linear}.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-HUofsb-Jt5cK{animation:mdc-checkbox-unchecked-checked-checkmark-path .18s linear 0s;transition:none}.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-SJnn3d{animation:mdc-checkbox-unchecked-indeterminate-mixedmark 90ms linear 0s;transition:none}.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-HUofsb-Jt5cK{animation:mdc-checkbox-checked-unchecked-checkmark-path 90ms linear 0s;transition:none}.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-A9y3zc .VfPpkd-HUofsb{animation:mdc-checkbox-checked-indeterminate-checkmark 90ms linear 0s;transition:none}.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-A9y3zc .VfPpkd-SJnn3d{animation:mdc-checkbox-checked-indeterminate-mixedmark 90ms linear 0s;transition:none}.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-barxie .VfPpkd-HUofsb{animation:mdc-checkbox-indeterminate-checked-checkmark .5s linear 0s;transition:none}.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-barxie .VfPpkd-SJnn3d{animation:mdc-checkbox-indeterminate-checked-mixedmark .5s linear 0s;transition:none}.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-SJnn3d{animation:mdc-checkbox-indeterminate-unchecked-mixedmark .3s linear 0s;transition:none}.VfPpkd-muHVFf-bMcfAe:checked~.VfPpkd-YQoJzd,.VfPpkd-muHVFf-bMcfAe:indeterminate~.VfPpkd-YQoJzd,.VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]~.VfPpkd-YQoJzd{transition:border-color 90ms 0ms cubic-bezier(0,0,.2,1),background-color 90ms 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-muHVFf-bMcfAe:checked~.VfPpkd-YQoJzd .VfPpkd-HUofsb-Jt5cK,.VfPpkd-muHVFf-bMcfAe:indeterminate~.VfPpkd-YQoJzd .VfPpkd-HUofsb-Jt5cK,.VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]~.VfPpkd-YQoJzd .VfPpkd-HUofsb-Jt5cK{stroke-dashoffset:0}.VfPpkd-muHVFf-bMcfAe{position:absolute;margin:0;padding:0;opacity:0;cursor:inherit}.VfPpkd-muHVFf-bMcfAe:disabled{cursor:default;pointer-events:none}.VfPpkd-MPu53c-OWXEXe-dgl2Hf{margin:4px;margin:calc((var(--mdc-checkbox-state-layer-size, 48px) - var(--mdc-checkbox-state-layer-size, 40px))/2)}.VfPpkd-MPu53c-OWXEXe-dgl2Hf .VfPpkd-muHVFf-bMcfAe{top:-4px;top:calc((var(--mdc-checkbox-state-layer-size, 40px) - var(--mdc-checkbox-state-layer-size, 48px))/2);right:-4px;right:calc((var(--mdc-checkbox-state-layer-size, 40px) - var(--mdc-checkbox-state-layer-size, 48px))/2);left:-4px;left:calc((var(--mdc-checkbox-state-layer-size, 40px) - var(--mdc-checkbox-state-layer-size, 48px))/2);width:48px;width:var(--mdc-checkbox-state-layer-size,48px);height:48px;height:var(--mdc-checkbox-state-layer-size,48px)}.VfPpkd-muHVFf-bMcfAe:checked~.VfPpkd-YQoJzd .VfPpkd-HUofsb{transition:opacity .18s 0ms cubic-bezier(0,0,.2,1),transform .18s 0ms cubic-bezier(0,0,.2,1);opacity:1}.VfPpkd-muHVFf-bMcfAe:checked~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{transform:scaleX(1) rotate(-45deg)}.VfPpkd-muHVFf-bMcfAe:indeterminate~.VfPpkd-YQoJzd .VfPpkd-HUofsb,.VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]~.VfPpkd-YQoJzd .VfPpkd-HUofsb{transform:rotate(45deg);opacity:0;transition:opacity 90ms 0ms cubic-bezier(.4,0,.6,1),transform 90ms 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-muHVFf-bMcfAe:indeterminate~.VfPpkd-YQoJzd .VfPpkd-SJnn3d,.VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{transform:scaleX(1) rotate(0deg);opacity:1}.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-YQoJzd,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-HUofsb,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-HUofsb-Jt5cK,.VfPpkd-MPu53c.VfPpkd-MPu53c-OWXEXe-mWPk3d .VfPpkd-SJnn3d{transition:none}.VfPpkd-MPu53c{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-MPu53c .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c .VfPpkd-OYHm6b::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-MPu53c .VfPpkd-OYHm6b::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-MPu53c .VfPpkd-OYHm6b::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-OYHm6b::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-OYHm6b::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-OYHm6b::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-MPu53c .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c .VfPpkd-OYHm6b::after{top:0;left:0;width:100%;height:100%}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0);width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-MPu53c.VfPpkd-ksKsZd-mWPk3d .VfPpkd-OYHm6b::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-MPu53c{z-index:0}.VfPpkd-MPu53c .VfPpkd-OYHm6b::before,.VfPpkd-MPu53c .VfPpkd-OYHm6b::after{z-index:-1;z-index:var(--mdc-ripple-z-index,-1)}.VfPpkd-OYHm6b{position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:GrayText;border-color:var(--mdc-checkbox-disabled-unselected-icon-color,GrayText);background-color:transparent}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:checked~.VfPpkd-YQoJzd,.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate~.VfPpkd-YQoJzd,.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true][disabled]~.VfPpkd-YQoJzd{border-color:GrayText;background-color:GrayText;background-color:var(--mdc-checkbox-disabled-selected-icon-color,GrayText)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:ButtonText;color:var(--mdc-checkbox-selected-checkmark-color,ButtonText)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:ButtonText;border-color:var(--mdc-checkbox-selected-checkmark-color,ButtonText)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:ButtonFace;color:var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace)}.VfPpkd-MPu53c .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:ButtonFace;border-color:var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace)}}.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgba(60,64,67,.38);border-color:var(--mdc-checkbox-disabled-unselected-icon-color,rgba(60,64,67,.38));background-color:transparent}.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:checked~.VfPpkd-YQoJzd,.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate~.VfPpkd-YQoJzd,.Ne8lhe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true][disabled]~.VfPpkd-YQoJzd{border-color:transparent;background-color:rgba(60,64,67,.38);background-color:var(--mdc-checkbox-disabled-selected-icon-color,rgba(60,64,67,.38))}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:#fff;color:var(--mdc-checkbox-selected-checkmark-color,#fff)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:#fff;border-color:var(--mdc-checkbox-selected-checkmark-color,#fff)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:#fff;color:var(--mdc-checkbox-disabled-selected-checkmark-color,#fff)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:#fff;border-color:var(--mdc-checkbox-disabled-selected-checkmark-color,#fff)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#5f6368;border-color:var(--mdc-checkbox-unselected-icon-color,#5f6368);background-color:transparent}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ne8lhe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#1a73e8;border-color:var(--mdc-checkbox-selected-icon-color,#1a73e8);background-color:#1a73e8;background-color:var(--mdc-checkbox-selected-icon-color,#1a73e8)}@keyframes mdc-checkbox-fade-in-background-FF5F6368FF1A73E800000000FF1A73E8{0%{border-color:#5f6368;border-color:var(--mdc-checkbox-unselected-icon-color,#5f6368);background-color:transparent}50%{border-color:#1a73e8;border-color:var(--mdc-checkbox-selected-icon-color,#1a73e8);background-color:#1a73e8;background-color:var(--mdc-checkbox-selected-icon-color,#1a73e8)}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FF1A73E800000000FF1A73E8{0%,80%{border-color:#1a73e8;border-color:var(--mdc-checkbox-selected-icon-color,#1a73e8);background-color:#1a73e8;background-color:var(--mdc-checkbox-selected-icon-color,#1a73e8)}100%{border-color:#5f6368;border-color:var(--mdc-checkbox-unselected-icon-color,#5f6368);background-color:transparent}}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FF1A73E800000000FF1A73E8}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FF1A73E800000000FF1A73E8}.Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#202124;border-color:var(--mdc-checkbox-unselected-hover-icon-color,#202124);background-color:transparent}.Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ne8lhe:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#174ea6;border-color:var(--mdc-checkbox-selected-hover-icon-color,#174ea6);background-color:#174ea6;background-color:var(--mdc-checkbox-selected-hover-icon-color,#174ea6)}.Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6}.Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6}.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#202124;border-color:var(--mdc-checkbox-unselected-focus-icon-color,#202124);background-color:transparent}.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#174ea6;border-color:var(--mdc-checkbox-selected-focus-icon-color,#174ea6);background-color:#174ea6;background-color:var(--mdc-checkbox-selected-focus-icon-color,#174ea6)}.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6}.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6}.Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#202124;border-color:var(--mdc-checkbox-unselected-pressed-icon-color,#202124);background-color:transparent}.Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ne8lhe:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#174ea6;border-color:var(--mdc-checkbox-selected-pressed-icon-color,#174ea6);background-color:#174ea6;background-color:var(--mdc-checkbox-selected-pressed-icon-color,#174ea6)}@keyframes mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6{0%{border-color:#202124;border-color:var(--mdc-checkbox-unselected-pressed-icon-color,#202124);background-color:transparent}50%{border-color:#174ea6;border-color:var(--mdc-checkbox-selected-pressed-icon-color,#174ea6);background-color:#174ea6;background-color:var(--mdc-checkbox-selected-pressed-icon-color,#174ea6)}}@keyframes mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6{0%,80%{border-color:#174ea6;border-color:var(--mdc-checkbox-selected-pressed-icon-color,#174ea6);background-color:#174ea6;background-color:var(--mdc-checkbox-selected-pressed-icon-color,#174ea6)}100%{border-color:#202124;border-color:var(--mdc-checkbox-unselected-pressed-icon-color,#202124);background-color:transparent}}.Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6}.Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ne8lhe:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6}.Ne8lhe .VfPpkd-OYHm6b::before,.Ne8lhe .VfPpkd-OYHm6b::after{background-color:#3c4043;background-color:var(--mdc-checkbox-unselected-hover-state-layer-color,#3c4043)}.Ne8lhe:hover .VfPpkd-OYHm6b::before,.Ne8lhe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before{opacity:.04;opacity:var(--mdc-checkbox-unselected-hover-state-layer-opacity,.04)}.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before,.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-checkbox-unselected-focus-state-layer-opacity,.12)}.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after{transition:opacity .15s linear}.Ne8lhe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-checkbox-unselected-pressed-state-layer-opacity,.1)}.Ne8lhe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-checkbox-unselected-pressed-state-layer-opacity,0.1)}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:#1a73e8;background-color:var(--mdc-checkbox-selected-hover-state-layer-color,#1a73e8)}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:hover .VfPpkd-OYHm6b::before,.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before{opacity:.04;opacity:var(--mdc-checkbox-selected-hover-state-layer-opacity,.04)}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before,.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-checkbox-selected-focus-state-layer-opacity,.12)}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after{transition:opacity .15s linear}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-checkbox-selected-pressed-state-layer-opacity,.1)}.Ne8lhe.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-checkbox-selected-pressed-state-layer-opacity,0.1)}.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.Ne8lhe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:#1a73e8;background-color:var(--mdc-checkbox-selected-hover-state-layer-color,#1a73e8)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:GrayText;border-color:var(--mdc-checkbox-disabled-unselected-icon-color,GrayText);background-color:transparent}.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:checked~.VfPpkd-YQoJzd,.Ne8lhe .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate~.VfPpkd-YQoJzd,.Ne8lhe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true][disabled]~.VfPpkd-YQoJzd{border-color:GrayText;background-color:GrayText;background-color:var(--mdc-checkbox-disabled-selected-icon-color,GrayText)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:ButtonText;color:var(--mdc-checkbox-selected-checkmark-color,ButtonText)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:ButtonText;border-color:var(--mdc-checkbox-selected-checkmark-color,ButtonText)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:ButtonFace;color:var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace)}.Ne8lhe .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:ButtonFace;border-color:var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace)}}.az2ine{will-change:unset}.VfPpkd-GCYh9b{padding:10px}.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgba(0,0,0,.54)}.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:#018786;border-color:var(--mdc-theme-secondary,#018786)}.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:#018786;border-color:var(--mdc-theme-secondary,#018786)}.VfPpkd-GCYh9b [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:disabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgba(0,0,0,.38)}.VfPpkd-GCYh9b [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:disabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgba(0,0,0,.38)}.VfPpkd-GCYh9b [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgba(0,0,0,.38)}.VfPpkd-GCYh9b .VfPpkd-RsCWK::before{background-color:#018786;background-color:var(--mdc-theme-secondary,#018786)}.VfPpkd-GCYh9b .VfPpkd-RsCWK::before{top:-10px;left:-10px;width:40px;height:40px}.VfPpkd-GCYh9b .VfPpkd-gBXA9-bMcfAe{top:0;right:0;left:0;width:40px;height:40px}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me .VfPpkd-gBXA9-bMcfAe:disabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:GrayText}.VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me .VfPpkd-gBXA9-bMcfAe:disabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:GrayText}.VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.VfPpkd-GCYh9b.VfPpkd-GCYh9b-OWXEXe-OWB6Me .VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:GrayText}}.VfPpkd-GCYh9b{display:inline-block;position:relative;-moz-box-flex:0;flex:0 0 auto;-moz-box-sizing:content-box;box-sizing:content-box;width:20px;height:20px;cursor:pointer;will-change:opacity,transform,border-color,color}.VfPpkd-GCYh9b[hidden]{display:none}.VfPpkd-RsCWK{display:inline-block;position:relative;-moz-box-sizing:border-box;box-sizing:border-box;width:20px;height:20px}.VfPpkd-RsCWK::before{position:absolute;transform:scale(0,0);border-radius:50%;opacity:0;pointer-events:none;content:"";transition:opacity .12s 0ms cubic-bezier(.4,0,.6,1),transform .12s 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-wVo5xe-LkdAo{position:absolute;top:0;left:0;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;border-width:2px;border-style:solid;border-radius:50%;transition:border-color .12s 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-Z5TpLc-LkdAo{position:absolute;top:0;left:0;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;transform:scale(0,0);border-width:10px;border-style:solid;border-radius:50%;transition:transform .12s 0ms cubic-bezier(.4,0,.6,1),border-color .12s 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-gBXA9-bMcfAe{position:absolute;margin:0;padding:0;opacity:0;cursor:inherit;z-index:1}.VfPpkd-GCYh9b-OWXEXe-dgl2Hf{margin-top:4px;margin-bottom:4px;margin-right:4px;margin-left:4px}.VfPpkd-GCYh9b-OWXEXe-dgl2Hf .VfPpkd-gBXA9-bMcfAe{top:-4px;right:-4px;left:-4px;width:48px;height:48px}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec,.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec{pointer-events:none;border:2px solid transparent;border-radius:6px;-moz-box-sizing:content-box;box-sizing:content-box;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:100%;width:100%}@media screen and (forced-colors:active){.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec,.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec{border-color:CanvasText}}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec::after,.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec::after{content:"";border:2px solid transparent;border-radius:8px;display:block;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-r6xRoe-LhBDec::after,.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-r6xRoe-LhBDec::after{border-color:CanvasText}}.VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK,.VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK{transition:opacity .12s 0ms cubic-bezier(0,0,.2,1),transform .12s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{transition:border-color .12s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{transition:transform .12s 0ms cubic-bezier(0,0,.2,1),border-color .12s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-GCYh9b-OWXEXe-OWB6Me{cursor:default;pointer-events:none}.VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{transform:scale(.5);transition:transform .12s 0ms cubic-bezier(0,0,.2,1),border-color .12s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK,[aria-disabled=true] .VfPpkd-gBXA9-bMcfAe+.VfPpkd-RsCWK{cursor:default}.VfPpkd-gBXA9-bMcfAe:focus+.VfPpkd-RsCWK::before{transform:scale(1);opacity:.12;transition:opacity .12s 0ms cubic-bezier(0,0,.2,1),transform .12s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-GCYh9b{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before,.VfPpkd-GCYh9b .VfPpkd-eHTEvd::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-GCYh9b .VfPpkd-eHTEvd::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-eHTEvd::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-eHTEvd::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-eHTEvd::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before,.VfPpkd-GCYh9b .VfPpkd-eHTEvd::after{top:0;left:0;width:100%;height:100%}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::before,.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0);width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-eHTEvd::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-GCYh9b .VfPpkd-eHTEvd::before,.VfPpkd-GCYh9b .VfPpkd-eHTEvd::after{background-color:#018786;background-color:var(--mdc-ripple-color,var(--mdc-theme-secondary,#018786))}.VfPpkd-GCYh9b:hover .VfPpkd-eHTEvd::before,.VfPpkd-GCYh9b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-eHTEvd::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-eHTEvd::after{transition:opacity .15s linear}.VfPpkd-GCYh9b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-eHTEvd::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-RsCWK::before,.VfPpkd-GCYh9b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-RsCWK::before{content:none}.VfPpkd-eHTEvd{position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}.kDzhGf{z-index:0}.kDzhGf .VfPpkd-eHTEvd::before,.kDzhGf .VfPpkd-eHTEvd::after{z-index:-1}.kDzhGf .VfPpkd-eHTEvd::before,.kDzhGf .VfPpkd-eHTEvd::after{background-color:rgb(26,115,232);background-color:var(--gm-radio-state-color,rgb(26,115,232))}.kDzhGf:hover .VfPpkd-eHTEvd::before,.kDzhGf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-eHTEvd::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-eHTEvd::after{transition:opacity .15s linear}.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-eHTEvd::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before,.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::after{background-color:rgb(60,64,67);background-color:var(--gm-radio-state-color,rgb(60,64,67))}.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before,.kDzhGf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before,.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::after{transition:opacity .15s linear}.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.kDzhGf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(95,99,104);border-color:var(--gm-radio-stroke-color--unchecked,rgb(95,99,104))}.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(26,115,232);border-color:var(--gm-radio-stroke-color--checked,rgb(26,115,232))}.kDzhGf .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(26,115,232);border-color:var(--gm-radio-ink-color,rgb(26,115,232))}.kDzhGf [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf .VfPpkd-gBXA9-bMcfAe:disabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgba(60,64,67,.38);border-color:var(--gm-radio-disabled-stroke-color--unchecked,rgba(60,64,67,.38))}.kDzhGf [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf .VfPpkd-gBXA9-bMcfAe:disabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgba(60,64,67,.38);border-color:var(--gm-radio-disabled-stroke-color--checked,rgba(60,64,67,.38))}.kDzhGf [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.kDzhGf .VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgba(60,64,67,.38);border-color:var(--gm-radio-disabled-ink-color,rgba(60,64,67,.38))}.kDzhGf .VfPpkd-RsCWK::before{background-color:rgb(26,115,232);background-color:var(--gm-radio-state-color,rgb(26,115,232))}.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf:active .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(32,33,36);border-color:var(--gm-radio-stroke-color--unchecked-stateful,rgb(32,33,36))}.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.kDzhGf:active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(23,78,166);border-color:var(--gm-radio-stroke-color--checked-stateful,rgb(23,78,166))}.kDzhGf:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.kDzhGf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.kDzhGf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.kDzhGf:active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(23,78,166);border-color:var(--gm-radio-ink-color--stateful,rgb(23,78,166))}.wHsUjf{will-change:unset}.VfPpkd-StrnGf-rymPhb{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);line-height:1.5rem;margin:0;padding:8px 0;list-style-type:none;color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87))}.VfPpkd-StrnGf-rymPhb:focus{outline:none}.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgba(0,0,0,.54);color:var(--mdc-theme-text-secondary-on-background,rgba(0,0,0,.54))}.VfPpkd-StrnGf-rymPhb-f7MjDc{background-color:transparent}.VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-icon-on-background,rgba(0,0,0,.38))}.VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38))}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc{padding-top:4px;padding-bottom:4px;font-size:.812rem}.VfPpkd-StrnGf-rymPhb-Tkg0ld{display:block}.VfPpkd-StrnGf-rymPhb-ibnC6b{display:-moz-box;display:flex;position:relative;-moz-box-align:center;align-items:center;-moz-box-pack:start;justify-content:flex-start;overflow:hidden;padding:0;padding-left:16px;padding-right:16px;height:48px}.VfPpkd-StrnGf-rymPhb-ibnC6b:focus{outline:none}.VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{border-color:CanvasText}}.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:3px double transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{border-color:CanvasText}}[dir=rtl] .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:72px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:0;padding-right:16px;height:72px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:20px;height:20px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-f7MjDc{flex-shrink:0;-moz-box-align:center;align-items:center;-moz-box-pack:center;justify-content:center;fill:currentColor;object-fit:cover;margin-left:0;margin-right:32px;width:24px;height:24px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:32px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:32px;width:24px;height:24px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:32px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:40px;height:40px;border-radius:50%}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:40px;height:40px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:56px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:100px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{display:-moz-inline-box;display:inline-flex}.VfPpkd-StrnGf-rymPhb-IhFlZd{margin-left:auto;margin-right:0}.VfPpkd-StrnGf-rymPhb-IhFlZd:not(.HzV7m-fuEl3d){-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit)}.VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl] .VfPpkd-StrnGf-rymPhb-IhFlZd,[dir=rtl] .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-IhFlZd{margin-left:0;margin-right:auto}.VfPpkd-StrnGf-rymPhb-b9t22c{text-overflow:ellipsis;white-space:nowrap;overflow:hidden}.VfPpkd-StrnGf-rymPhb-b9t22c[for]{pointer-events:none}.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden;display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:24px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit);text-overflow:ellipsis;white-space:nowrap;overflow:hidden;display:block;margin-top:0;line-height:normal}.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{font-size:inherit}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b{height:40px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc .VfPpkd-StrnGf-rymPhb-b9t22c{align-self:flex-start}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc .VfPpkd-StrnGf-rymPhb-ibnC6b{height:64px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{height:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{align-self:flex-start;margin-top:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b{height:60px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:36px;height:36px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b{cursor:pointer}a.VfPpkd-StrnGf-rymPhb-ibnC6b{color:inherit;text-decoration:none}.VfPpkd-StrnGf-rymPhb-clz4Ic{height:0;margin:0;border:none;border-bottom-width:1px;border-bottom-style:solid}.VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(0,0,0,.12)}.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd,.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe,.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd,.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:88px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:88px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:88px;margin-right:0;width:calc(100% - 104px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:88px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:116px;margin-right:0;width:calc(100% - 116px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:116px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:116px;margin-right:0;width:calc(100% - 132px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:116px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:0;margin-right:0;width:100%}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:0;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:0}.VfPpkd-StrnGf-rymPhb-JNdkSc .VfPpkd-StrnGf-rymPhb{padding:0}.VfPpkd-StrnGf-rymPhb-oT7voc{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);margin:.75rem 16px}.VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87))}.VfPpkd-rymPhb-L8ivfd-fmcmS{color:rgba(0,0,0,.54);color:var(--mdc-theme-text-secondary-on-background,rgba(0,0,0,.54))}.VfPpkd-rymPhb-bC5pod-fmcmS{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38))}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{background-color:transparent}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-icon-on-background,rgba(0,0,0,.38))}.VfPpkd-rymPhb-JMEf7e{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38))}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-StrnGf-rymPhb-oT7voc{color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87))}.VfPpkd-rymPhb-clz4Ic::after{border-bottom-color:white}.VfPpkd-rymPhb{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);line-height:1.5rem}.VfPpkd-rymPhb-fpDzbe-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit)}.VfPpkd-rymPhb-L8ivfd-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit)}.VfPpkd-rymPhb-bC5pod-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-overline-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-overline-font-size,.75rem);line-height:2rem;line-height:var(--mdc-typography-overline-line-height,2rem);font-weight:500;font-weight:var(--mdc-typography-overline-font-weight,500);letter-spacing:.1666666667em;letter-spacing:var(--mdc-typography-overline-letter-spacing,.1666666667em);text-decoration:none;-moz-text-decoration:var(--mdc-typography-overline-text-decoration,none);text-decoration:var(--mdc-typography-overline-text-decoration,none);text-transform:uppercase;text-transform:var(--mdc-typography-overline-text-transform,uppercase)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{width:24px;height:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb{width:56px;height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb{width:100px;height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb{width:36px;height:20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{width:24px;height:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e{width:36px;height:20px}.VfPpkd-rymPhb-oT7voc{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit)}.VfPpkd-rymPhb-clz4Ic{background-color:rgba(0,0,0,.12)}.VfPpkd-rymPhb-clz4Ic{height:1px}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-rymPhb-clz4Ic::after{content:"";display:block;border-bottom-width:1px;border-bottom-style:solid}}.VfPpkd-rymPhb{margin:0;padding:8px 0;list-style-type:none}.VfPpkd-rymPhb:focus{outline:none}.VfPpkd-rymPhb-Tkg0ld{display:block}.VfPpkd-rymPhb-ibnC6b{display:-moz-box;display:flex;position:relative;-moz-box-align:center;align-items:center;-moz-box-pack:start;justify-content:flex-start;overflow:hidden;padding:0;-moz-box-align:stretch;align-items:stretch;cursor:pointer}.VfPpkd-rymPhb-ibnC6b:focus{outline:none}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:48px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:64px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb{height:88px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc .VfPpkd-rymPhb-KkROqb{align-self:center;margin-top:0}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e{align-self:center;margin-top:0}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me,.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-tPcied-hXIJHe{cursor:auto}.VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{border-color:CanvasText}}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:3px double transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{border-color:CanvasText}}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:focus::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:3px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:focus::before{border-color:CanvasText}}a.VfPpkd-rymPhb-ibnC6b{color:inherit;text-decoration:none}.VfPpkd-rymPhb-KkROqb{fill:currentColor;flex-shrink:0;pointer-events:none}.VfPpkd-rymPhb-JMEf7e{flex-shrink:0;pointer-events:none}.VfPpkd-rymPhb-Gtdoyb{text-overflow:ellipsis;white-space:nowrap;overflow:hidden;align-self:center;-moz-box-flex:1;flex:1;pointer-events:none}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-Gtdoyb{align-self:stretch}.VfPpkd-rymPhb-Gtdoyb[for]{pointer-events:none}.VfPpkd-rymPhb-fpDzbe-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-L8ivfd-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden;display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-L8ivfd-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS{white-space:normal;line-height:20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj .VfPpkd-rymPhb-L8ivfd-fmcmS{white-space:nowrap;line-height:auto}.VfPpkd-rymPhb-bC5pod-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:24px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb{border-radius:50%}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:32px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:32px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb{margin-left:0;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:24px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:24px;margin-right:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:24px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:24px;margin-right:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{align-self:flex-start;margin-top:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{margin-left:28px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:28px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e{margin-left:24px;margin-right:8px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:8px;margin-right:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e{margin-left:24px;margin-right:8px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:8px;margin-right:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b{padding-left:16px;padding-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-rymPhb-JNdkSc .VfPpkd-StrnGf-rymPhb{padding:0}.VfPpkd-rymPhb-oT7voc{margin:.75rem 16px}.VfPpkd-rymPhb-clz4Ic{padding:0;background-clip:content-box}.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe{padding-left:16px;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl]{padding-left:auto;padding-right:16px}.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe{padding-left:auto;padding-right:16px}[dir=rtl] .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl]{padding-left:16px;padding-right:auto}.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl]{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-clz4Ic,.VfPpkd-rymPhb-clz4Ic[dir=rtl]{padding:0}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::before{transform:scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:0;left:0;transform:scale(0);transform-origin:center center}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-StrnGf-rymPhb-pZXsl::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-StrnGf-rymPhb-pZXsl::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::before{transform:scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{top:0;left:0;transform:scale(0);transform-origin:center center}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-rymPhb-pZXsl::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-rymPhb-pZXsl::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-activated-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-activated-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.08;opacity:var(--mdc-ripple-selected-opacity,.08)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-hover-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-focus-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:.08;opacity:var(--mdc-ripple-selected-opacity,.08)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-hover-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-focus-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl{position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-StrnGf-rymPhb-pZXsl::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-StrnGf-rymPhb-pZXsl::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-rymPhb-pZXsl::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-rymPhb-pZXsl::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-pZXsl,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-pZXsl{position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::before{transform:scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{top:0;left:0;transform:scale(0);transform-origin:center center}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-rymPhb-pZXsl::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-rymPhb-pZXsl::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-activated-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:.08;opacity:var(--mdc-ripple-selected-opacity,.08)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-hover-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-focus-opacity,.2)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl{position:relative;outline:none;overflow:hidden;position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}.P2Hi5d,.mkMxfe,.OBi8lb,.P9QRxe,.vqjb4e,.y8Rdrf,.DMZ54e{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:#000;color:var(--mdc-theme-on-surface,#000)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-IhFlZd,.mkMxfe .VfPpkd-StrnGf-rymPhb-IhFlZd,.OBi8lb .VfPpkd-StrnGf-rymPhb-IhFlZd,.P9QRxe .VfPpkd-StrnGf-rymPhb-IhFlZd,.vqjb4e .VfPpkd-StrnGf-rymPhb-IhFlZd,.y8Rdrf .VfPpkd-StrnGf-rymPhb-IhFlZd,.DMZ54e .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(95,99,104)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(60,64,67)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#000;color:var(--mdc-theme-on-surface,#000)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#000;color:var(--mdc-theme-on-surface,#000)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:24px;padding-right:16px}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:24px;margin-right:0;width:calc(100% - 24px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:24px;margin-right:0;width:calc(100% - 40px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:24px;margin-right:0;width:calc(100% - 24px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:24px;margin-right:0;width:calc(100% - 40px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:24px}.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:56px;margin-right:0;width:calc(100% - 56px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:56px}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:56px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:56px}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.r6B9Fd{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400}.r6B9Fd .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(60,64,67)}.r6B9Fd .VfPpkd-rymPhb-L8ivfd-fmcmS,.r6B9Fd .VfPpkd-rymPhb-bC5pod-fmcmS,.r6B9Fd .VfPpkd-rymPhb-JMEf7e{color:rgb(95,99,104)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:rgb(60,64,67)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:rgb(60,64,67)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:0}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media screen and (forced-colors:active){.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:GrayText}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:1}}.uTZ9Lb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.FvXOfd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.QrsYgb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.gfwIBd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:center;margin-top:0}.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:72px}.UbEQCe.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .UbEQCe.VfPpkd-rymPhb-ibnC6b,.UbEQCe.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.UbEQCe .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .UbEQCe .VfPpkd-rymPhb-KkROqb,.UbEQCe .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.rKASPc.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .rKASPc.VfPpkd-rymPhb-ibnC6b,.rKASPc.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.rKASPc .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:8px}[dir=rtl] .rKASPc .VfPpkd-rymPhb-KkROqb,.rKASPc .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:8px;margin-right:8px}.rKASPc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:8px}.U5k4Fd.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .U5k4Fd.VfPpkd-rymPhb-ibnC6b,.U5k4Fd.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.U5k4Fd .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:8px}[dir=rtl] .U5k4Fd .VfPpkd-rymPhb-KkROqb,.U5k4Fd .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:8px;margin-right:8px}.U5k4Fd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:8px}.ifEyr.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .ifEyr.VfPpkd-rymPhb-ibnC6b,.ifEyr.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.ifEyr .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:8px}[dir=rtl] .ifEyr .VfPpkd-rymPhb-KkROqb,.ifEyr .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:8px;margin-right:8px}.ifEyr.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{align-self:flex-start;margin-top:8px}.SNowt.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .SNowt.VfPpkd-rymPhb-ibnC6b,.SNowt.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.SNowt .VfPpkd-rymPhb-JMEf7e{margin-left:8px;margin-right:16px}[dir=rtl] .SNowt .VfPpkd-rymPhb-JMEf7e,.SNowt .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:8px}.tfmWAf.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .tfmWAf.VfPpkd-rymPhb-ibnC6b,.tfmWAf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.tfmWAf .VfPpkd-rymPhb-JMEf7e{margin-left:8px;margin-right:16px}[dir=rtl] .tfmWAf .VfPpkd-rymPhb-JMEf7e,.tfmWAf .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:8px}.axtYbd.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .axtYbd.VfPpkd-rymPhb-ibnC6b,.axtYbd.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.axtYbd .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:24px}[dir=rtl] .axtYbd .VfPpkd-rymPhb-JMEf7e,.axtYbd .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:24px;margin-right:16px}.aopLEb.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .aopLEb.VfPpkd-rymPhb-ibnC6b,.aopLEb.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.aopLEb .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:24px}[dir=rtl] .aopLEb .VfPpkd-rymPhb-JMEf7e,.aopLEb .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:24px;margin-right:16px}.zlqiud.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .zlqiud.VfPpkd-rymPhb-ibnC6b,.zlqiud.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.zlqiud .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:24px}[dir=rtl] .zlqiud .VfPpkd-rymPhb-JMEf7e,.zlqiud .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:24px;margin-right:16px}.isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe{padding-left:24px;padding-right:auto}[dir=rtl] .isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl]{padding-left:auto;padding-right:24px}.MCs1Pd{padding-left:24px;padding-right:24px}[dir=rtl] .MCs1Pd,.MCs1Pd[dir=rtl]{padding-left:24px;padding-right:24px}.e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe{padding-left:auto;padding-right:24px}[dir=rtl] .e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl]{padding-left:24px;padding-right:auto}[dir=rtl] .e6pQl,.e6pQl[dir=rtl]{padding:0}.VfPpkd-xl07Ob-XxIAqe{display:none;position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;margin:0;padding:0;transform:scale(1);transform-origin:top left;opacity:0;overflow:auto;will-change:transform,opacity;box-shadow:0 5px 5px -3px rgba(0,0,0,.2),0 8px 10px 1px rgba(0,0,0,.14),0 3px 14px 2px rgba(0,0,0,.12);transform-origin-left:top left;transform-origin-right:top right}.VfPpkd-xl07Ob-XxIAqe:focus{outline:none}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-FNFY6c{display:inline-block;transform:scale(.8);opacity:0}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-FNFY6c{display:inline-block;transform:scale(1);opacity:1}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-xTMeO{display:inline-block;opacity:0}[dir=rtl] .VfPpkd-xl07Ob-XxIAqe,.VfPpkd-xl07Ob-XxIAqe[dir=rtl]{transform-origin-left:top right;transform-origin-right:top left}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd{position:relative;overflow:visible}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL{position:fixed}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-tsQazb{width:100%}.VfPpkd-xl07Ob-XxIAqe{max-width:calc(100vw - 32px);max-width:var(--mdc-menu-max-width,calc(100vw - 32px));max-height:calc(100vh - 32px);max-height:var(--mdc-menu-max-height,calc(100vh - 32px));z-index:8;transition:opacity .03s linear,transform .12s cubic-bezier(0,0,.2,1),height .25s cubic-bezier(0,0,.2,1);background-color:#fff;background-color:var(--mdc-theme-surface,#fff);color:#000;color:var(--mdc-theme-on-surface,#000);border-radius:4px;border-radius:var(--mdc-shape-medium,4px)}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-xTMeO{transition:opacity 75ms linear}.VfPpkd-xl07Ob{min-width:112px;min-width:var(--mdc-menu-min-width,112px)}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-IhFlZd,.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgba(0,0,0,.87)}.VfPpkd-xl07Ob .VfPpkd-xl07Ob-ibnC6b-OWXEXe-eKm5Fc-FNFY6c .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04}.VfPpkd-xl07Ob .VfPpkd-xl07Ob-ibnC6b-OWXEXe-eKm5Fc-FNFY6c .VfPpkd-rymPhb-pZXsl::before{opacity:.04}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb{color:rgba(0,0,0,.87)}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb,.VfPpkd-xl07Ob .VfPpkd-rymPhb{position:relative}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb .VfPpkd-BFbNVe-bF1uUb,.VfPpkd-xl07Ob .VfPpkd-rymPhb .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb::before,.VfPpkd-xl07Ob .VfPpkd-rymPhb::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb::before,.VfPpkd-xl07Ob .VfPpkd-rymPhb::before{border-color:CanvasText}}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-clz4Ic{margin:8px 0}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-ibnC6b{-moz-user-select:none;user-select:none}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me{cursor:auto}.VfPpkd-xl07Ob a.VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-b9t22c,.VfPpkd-xl07Ob a.VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{pointer-events:none}.VfPpkd-qPzbhe-JNdkSc{padding:0;fill:currentColor}.VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:56px;padding-right:16px}[dir=rtl] .VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:56px}.VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c{left:16px;right:auto;display:none;position:absolute;top:50%;transform:translateY(-50%)}[dir=rtl] .VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c,.VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c[dir=rtl]{left:auto;right:16px}.VfPpkd-xl07Ob-ibnC6b-OWXEXe-gk6SMd .VfPpkd-qPzbhe-JNdkSc-Bz112c{display:inline}.O1htCb-H9tDt{display:-moz-inline-box;display:inline-flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;position:relative}.O1htCb-H9tDt[hidden]{display:none}@charset "UTF-8";.VfPpkd-O1htCb{display:-moz-inline-box;display:inline-flex;position:relative}.VfPpkd-O1htCb .VfPpkd-NLUYnc-V67aGc{top:50%;transform:translateY(-50%);pointer-events:none}.VfPpkd-O1htCb .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px}[dir=rtl] .VfPpkd-O1htCb .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-O1htCb .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-O1htCb .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:12px}[dir=rtl] .VfPpkd-O1htCb .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-O1htCb .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:12px;margin-right:0}.VfPpkd-O1htCb[hidden]{display:none}.VfPpkd-t08AT-Bz112c{display:-moz-inline-box;display:inline-flex;position:relative;align-self:center;-moz-box-align:center;align-items:center;-moz-box-pack:center;justify-content:center;flex-shrink:0;pointer-events:none}.VfPpkd-t08AT-Bz112c .VfPpkd-t08AT-Bz112c-auswjd,.VfPpkd-t08AT-Bz112c .VfPpkd-t08AT-Bz112c-mt1Mkb{position:absolute;top:0;left:0}.VfPpkd-t08AT-Bz112c .VfPpkd-t08AT-Bz112c-Bd00G{width:41.6666666667%;height:20.8333333333%}.VfPpkd-t08AT-Bz112c .VfPpkd-t08AT-Bz112c-mt1Mkb{opacity:1;transition:opacity 75ms linear 75ms}.VfPpkd-t08AT-Bz112c .VfPpkd-t08AT-Bz112c-auswjd{opacity:0;transition:opacity 75ms linear}.VfPpkd-O1htCb-OWXEXe-pXU01b .VfPpkd-t08AT-Bz112c .VfPpkd-t08AT-Bz112c-mt1Mkb{opacity:0;transition:opacity 49.5ms linear}.VfPpkd-O1htCb-OWXEXe-pXU01b .VfPpkd-t08AT-Bz112c .VfPpkd-t08AT-Bz112c-auswjd{opacity:1;transition:opacity .1005s linear 49.5ms}.VfPpkd-TkwUic{min-width:0;-moz-box-flex:1;flex:1 1 auto;position:relative;-moz-box-sizing:border-box;box-sizing:border-box;overflow:hidden;outline:none;cursor:pointer}.VfPpkd-uusGie-fmcmS-haAclf{display:-moz-box;display:flex;-moz-appearance:none;appearance:none;pointer-events:none;-moz-box-sizing:border-box;box-sizing:border-box;width:auto;min-width:0;-moz-box-flex:1;flex-grow:1;border:none;outline:none;padding:0;background-color:transparent;color:inherit}.VfPpkd-uusGie-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);text-overflow:ellipsis;white-space:nowrap;overflow:hidden;display:block;width:100%;text-align:left}[dir=rtl] .VfPpkd-uusGie-fmcmS,.VfPpkd-uusGie-fmcmS[dir=rtl]{text-align:right}.VfPpkd-O1htCb-OWXEXe-OWB6Me{cursor:default;pointer-events:none}.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:12px;padding-right:12px}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:12px;padding-right:12px}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-YPmvEd::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}}@media screen and (-ms-high-contrast:active) and (forced-colors:active),screen and (forced-colors:active) and (forced-colors:active){.VfPpkd-YPmvEd::before{border-color:CanvasText}}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-cTi5dd,.VfPpkd-YPmvEd .VfPpkd-rymPhb .VfPpkd-cTi5dd{margin-left:0;margin-right:0}[dir=rtl] .VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-cTi5dd,[dir=rtl] .VfPpkd-YPmvEd .VfPpkd-rymPhb .VfPpkd-cTi5dd,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-cTi5dd[dir=rtl],.VfPpkd-YPmvEd .VfPpkd-rymPhb .VfPpkd-cTi5dd[dir=rtl]{margin-left:0;margin-right:0}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.VfPpkd-YPmvEd .VfPpkd-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.VfPpkd-YPmvEd .VfPpkd-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-YPmvEd .VfPpkd-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-YPmvEd .VfPpkd-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-YPmvEd .VfPpkd-rymPhb-KkROqb{display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center}.VfPpkd-OkbHre{padding-left:16px;padding-right:16px}[dir=rtl] .VfPpkd-OkbHre,.VfPpkd-OkbHre[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-aJasdd-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:48px}.VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:64px}.VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{margin-top:20px}.VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:36px;content:"";vertical-align:0}.VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc{padding-left:0;padding-right:12px}.VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc.VfPpkd-rymPhb-ibnC6b,.VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc .VfPpkd-rymPhb-KkROqb{margin-left:12px;margin-right:0}[dir=rtl] .VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc .VfPpkd-rymPhb-KkROqb,.VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:0;margin-right:12px}.VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc .VfPpkd-rymPhb-KkROqb{width:36px;height:24px}[dir=rtl] .VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc,.VfPpkd-OkbHre-SfQLQb-M1Soyc-bN97Pc[dir=rtl]{padding-left:12px;padding-right:0}.VfPpkd-OkbHre-SfQLQb-r4m2rf.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-OkbHre-SfQLQb-r4m2rf.VfPpkd-rymPhb-ibnC6b,.VfPpkd-OkbHre-SfQLQb-r4m2rf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-OkbHre-SfQLQb-r4m2rf .VfPpkd-rymPhb-JMEf7e{margin-left:12px;margin-right:12px}[dir=rtl] .VfPpkd-OkbHre-SfQLQb-r4m2rf .VfPpkd-rymPhb-JMEf7e,.VfPpkd-OkbHre-SfQLQb-r4m2rf .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:12px;margin-right:12px}.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-xl07Ob-XxIAqe-OWXEXe-uxVfW-FNFY6c-uFfGwd{border-top-left-radius:0;border-top-right-radius:0}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-XpnDCe.VfPpkd-RWgCYc-ksKsZd::after{transform:scale(1,2);opacity:1}.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-TkwUic{height:56px;display:-moz-box;display:flex;-moz-box-align:baseline;align-items:baseline}.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-TkwUic::before{display:inline-block;width:0;height:40px;content:"";vertical-align:0}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS::before{content:"​"}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS-haAclf{height:100%;display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic::before{display:none}.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-TkwUic{border-top-left-radius:4px;border-top-left-radius:var(--mdc-shape-small,4px);border-top-right-radius:4px;border-top-right-radius:var(--mdc-shape-small,4px);border-bottom-right-radius:0;border-bottom-left-radius:0}.VfPpkd-O1htCb-OWXEXe-MFS4be:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-TkwUic{background-color:whitesmoke}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-TkwUic{background-color:#fafafa}.VfPpkd-O1htCb-OWXEXe-MFS4be:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(0,0,0,.42)}.VfPpkd-O1htCb-OWXEXe-MFS4be:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(0,0,0,.87)}.VfPpkd-O1htCb-OWXEXe-MFS4be:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:#6200ee;border-bottom-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(0,0,0,.06)}.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{max-width:calc(100% - 64px)}.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:calc(133.3333333333% - 85.3333333333px)}.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{left:16px;right:auto}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc,.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:16px}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc{left:48px;right:auto}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc,.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:48px}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc{max-width:calc(100% - 96px)}.VfPpkd-O1htCb-OWXEXe-MFS4be.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:calc(133.3333333333% - 128px)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:#b00020;border-bottom-color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:#b00020;border-bottom-color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:#b00020;border-bottom-color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-INsAgc{border:none}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic{display:-moz-box;display:flex;-moz-box-align:baseline;align-items:baseline;overflow:visible}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-uusGie-fmcmS-haAclf{display:-moz-box;display:flex;border:none;z-index:1;background-color:transparent}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-cTi5dd{z-index:2}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-xl07Ob-XxIAqe{margin-bottom:8px}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-xl07Ob-XxIAqe,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-xl07Ob-XxIAqe-OWXEXe-uxVfW-FNFY6c-uFfGwd{margin-bottom:0}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic{height:56px}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-select-outlined-56px .25s 1}@keyframes mdc-floating-label-shake-float-above-select-outlined-56px{0%{transform:translateX(0) translateY(-34.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(4%) translateY(-34.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(-4%) translateY(-34.75px) scale(.75)}100%{transform:translateX(0) translateY(-34.75px) scale(.75)}}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb{border-top-left-radius:4px;border-top-left-radius:var(--mdc-shape-small,4px);border-top-right-radius:0;border-bottom-right-radius:0;border-bottom-left-radius:4px;border-bottom-left-radius:var(--mdc-shape-small,4px)}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb[dir=rtl]{border-top-left-radius:0;border-top-right-radius:4px;border-top-right-radius:var(--mdc-shape-small,4px);border-bottom-right-radius:4px;border-bottom-right-radius:var(--mdc-shape-small,4px);border-bottom-left-radius:0}@supports (top:max(0%)){.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb{width:max(12px,var(--mdc-shape-small,4px))}}@supports (top:max(0%)){.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd{max-width:calc(100% - max(12px, var(--mdc-shape-small, 4px))*2)}}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-top-left-radius:0;border-top-right-radius:4px;border-top-right-radius:var(--mdc-shape-small,4px);border-bottom-right-radius:4px;border-bottom-right-radius:var(--mdc-shape-small,4px);border-bottom-left-radius:0}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe[dir=rtl]{border-top-left-radius:4px;border-top-left-radius:var(--mdc-shape-small,4px);border-top-right-radius:0;border-bottom-right-radius:0;border-bottom-left-radius:4px;border-bottom-left-radius:var(--mdc-shape-small,4px)}@supports (top:max(0%)){.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic{padding-left:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic[dir=rtl]{padding-left:0}@supports (top:max(0%)){[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic[dir=rtl]{padding-right:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}@supports (top:max(0%)){.VfPpkd-O1htCb-OWXEXe-INsAgc+.VfPpkd-O1htCb-W0vJo-fmcmS{margin-left:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc+.VfPpkd-O1htCb-W0vJo-fmcmS,.VfPpkd-O1htCb-OWXEXe-INsAgc+.VfPpkd-O1htCb-W0vJo-fmcmS[dir=rtl]{margin-left:0}@supports (top:max(0%)){[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc+.VfPpkd-O1htCb-W0vJo-fmcmS,.VfPpkd-O1htCb-OWXEXe-INsAgc+.VfPpkd-O1htCb-W0vJo-fmcmS[dir=rtl]{margin-right:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-TkwUic{background-color:transparent}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-TkwUic{background-color:transparent}.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(0,0,0,.38)}.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(0,0,0,.87)}.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:#6200ee;border-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(0,0,0,.06)}.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-width:2px}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic :not(.VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd) .VfPpkd-NSFCdd-Ra9xwd{max-width:calc(100% - 60px)}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-select-outlined .25s 1}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-37.25px) scale(1)}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:.75rem}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-34.75px) scale(.75)}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:1rem}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd{padding-top:1px}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS::before{content:"​"}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS-haAclf{height:100%;display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-TkwUic::before{display:none}.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc{line-height:1.15rem;left:4px;right:auto}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc,.VfPpkd-O1htCb-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:4px}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd{padding-top:2px}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:#b00020;border-color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:#b00020;border-color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:#b00020;border-color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc{left:36px;right:auto}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:36px}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-37.25px) translateX(-32px) scale(1)}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe[dir=rtl]{transform:translateY(-37.25px) translateX(32px) scale(1)}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:.75rem}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-34.75px) translateX(-32px) scale(.75)}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe[dir=rtl],.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe[dir=rtl]{transform:translateY(-34.75px) translateX(32px) scale(.75)}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:1rem}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-select-outlined-leading-icon-56px .25s 1}@keyframes mdc-floating-label-shake-float-above-select-outlined-leading-icon-56px{0%{transform:translateX(-32px) translateY(-34.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(calc(4% - 32px)) translateY(-34.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(calc(-4% - 32px)) translateY(-34.75px) scale(.75)}100%{transform:translateX(-32px) translateY(-34.75px) scale(.75)}}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU,.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c[dir=rtl] .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-select-outlined-leading-icon-56px .25s 1}@keyframes mdc-floating-label-shake-float-above-select-outlined-leading-icon-56px-rtl{0%{transform:translateX(32px) translateY(-34.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(calc(4% + 32px)) translateY(-34.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(calc(-4% + 32px)) translateY(-34.75px) scale(.75)}100%{transform:translateX(32px) translateY(-34.75px) scale(.75)}}.VfPpkd-O1htCb-OWXEXe-INsAgc.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-TkwUic :not(.VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd) .VfPpkd-NSFCdd-Ra9xwd{max-width:calc(100% - 96px)}.VfPpkd-TkwUic{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-TkwUic .VfPpkd-woaZLe::before,.VfPpkd-TkwUic .VfPpkd-woaZLe::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-TkwUic .VfPpkd-woaZLe::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-TkwUic .VfPpkd-woaZLe::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d .VfPpkd-woaZLe::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d .VfPpkd-woaZLe::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-woaZLe::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-woaZLe::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-woaZLe::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-TkwUic .VfPpkd-woaZLe::before,.VfPpkd-TkwUic .VfPpkd-woaZLe::after{top:-50%;left:-50%;width:200%;height:200%}.VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d .VfPpkd-woaZLe::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-TkwUic .VfPpkd-woaZLe::before,.VfPpkd-TkwUic .VfPpkd-woaZLe::after{background-color:rgba(0,0,0,.87);background-color:var(--mdc-ripple-color,rgba(0,0,0,.87))}.VfPpkd-TkwUic:hover .VfPpkd-woaZLe::before,.VfPpkd-TkwUic.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-woaZLe::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-woaZLe::before,.VfPpkd-TkwUic:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-woaZLe::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-TkwUic .VfPpkd-woaZLe{position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-YPmvEd .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-O1htCb-W0vJo-fmcmS{margin:0;margin-left:16px;margin-right:16px;-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit);display:block;margin-top:0;line-height:normal}[dir=rtl] .VfPpkd-O1htCb-W0vJo-fmcmS,.VfPpkd-O1htCb-W0vJo-fmcmS[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-O1htCb-W0vJo-fmcmS::before{display:inline-block;width:0;height:16px;content:"";vertical-align:0}.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{opacity:0;transition:opacity .18s cubic-bezier(.4,0,.2,1)}.VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb,.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb-zvnfze{opacity:1}.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-cTi5dd{display:inline-block;-moz-box-sizing:border-box;box-sizing:border-box;border:none;text-decoration:none;cursor:pointer;-moz-user-select:none;user-select:none;flex-shrink:0;align-self:center;background-color:transparent;fill:currentColor}.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-cTi5dd{margin-left:12px;margin-right:12px}[dir=rtl] .VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-cTi5dd,.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-cTi5dd[dir=rtl]{margin-left:12px;margin-right:12px}.VfPpkd-cTi5dd:not([tabindex]),.VfPpkd-cTi5dd[tabindex="-1"]{cursor:default;pointer-events:none}.VfPpkd-O1htCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-uusGie-fmcmS{color:rgba(0,0,0,.87)}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:rgba(0,0,0,.38)}.VfPpkd-O1htCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgba(0,0,0,.6)}.VfPpkd-O1htCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgba(98,0,238,.87)}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(0,0,0,.38)}.VfPpkd-O1htCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgba(0,0,0,.54)}.VfPpkd-O1htCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:#6200ee;fill:var(--mdc-theme-primary,#6200ee)}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-t08AT-Bz112c{fill:rgba(0,0,0,.38)}.VfPpkd-O1htCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me)+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgba(0,0,0,.6)}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgba(0,0,0,.38)}.VfPpkd-O1htCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-cTi5dd{color:rgba(0,0,0,.54)}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-cTi5dd{color:rgba(0,0,0,.38)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:GrayText}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-t08AT-Bz112c{fill:red}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:GrayText}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:GrayText}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:GrayText}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-cTi5dd,.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-OWB6Me+.VfPpkd-O1htCb-W0vJo-fmcmS{color:GrayText}}.VfPpkd-O1htCb .VfPpkd-TkwUic{padding-left:16px;padding-right:0}[dir=rtl] .VfPpkd-O1htCb .VfPpkd-TkwUic,.VfPpkd-O1htCb .VfPpkd-TkwUic[dir=rtl]{padding-left:0;padding-right:16px}.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-TkwUic{padding-left:0;padding-right:0}[dir=rtl] .VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-TkwUic,.VfPpkd-O1htCb.VfPpkd-O1htCb-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-TkwUic[dir=rtl]{padding-left:0;padding-right:0}.VfPpkd-O1htCb .VfPpkd-cTi5dd{width:24px;height:24px;font-size:24px}.VfPpkd-O1htCb .VfPpkd-t08AT-Bz112c{width:24px;height:24px}.VfPpkd-t08AT-Bz112c{margin-left:12px;margin-right:12px}[dir=rtl] .VfPpkd-t08AT-Bz112c,.VfPpkd-t08AT-Bz112c[dir=rtl]{margin-left:12px;margin-right:12px}.VfPpkd-TkwUic{width:200px}.VfPpkd-TkwUic .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-106%) scale(.75)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:#b00020;color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:#b00020;color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:#b00020;color:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:#b00020;fill:var(--mdc-theme-error,#b00020)}.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:#b00020;fill:var(--mdc-theme-error,#b00020)}.VfPpkd-uusGie-fmcmS-haAclf{height:28px}.s8kOBc{box-shadow:0 3px 5px -1px rgba(0,0,0,.2),0 6px 10px 0 rgba(0,0,0,.14),0 1px 18px 0 rgba(0,0,0,.12);font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400}.s8kOBc .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:rgb(60,64,67)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(95,99,104)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(60,64,67)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(60,64,67)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}.s8kOBc .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(60,64,67)}.s8kOBc .VfPpkd-rymPhb-L8ivfd-fmcmS,.s8kOBc .VfPpkd-rymPhb-bC5pod-fmcmS,.s8kOBc .VfPpkd-rymPhb-JMEf7e{color:rgb(95,99,104)}.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:rgb(60,64,67)}.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:rgb(60,64,67)}.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:0}.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.s8kOBc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media screen and (forced-colors:active){.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:GrayText}.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.s8kOBc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:1}}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(95,99,104)}.s8kOBc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.s8kOBc .VfPpkd-rymPhb .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.s8kOBc .VfPpkd-rymPhb .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:rgb(60,64,67)}.s8kOBc .VfPpkd-rymPhb-fpDzbe-fmcmS{letter-spacing:.00625em}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(252,232,230)}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(217,48,37);background-color:var(--mdc-ripple-color,rgb(217,48,37))}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(217,48,37);background-color:var(--mdc-ripple-color,rgb(217,48,37))}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{transition:opacity .15s linear}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.s8kOBc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-TkwUic{background-color:rgb(241,243,244)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-TkwUic{background-color:rgba(95,99,104,.04)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(95,99,104)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(32,33,36)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(25,103,210)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(95,99,104,.38)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(95,99,104)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(25,103,210)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(32,33,36)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(95,99,104,.38)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me)+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgb(95,99,104)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-OWB6Me+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgba(95,99,104,.38)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(197,34,31)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover.VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(165,14,14)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-uusGie-fmcmS{color:rgb(60,64,67)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:rgba(60,64,67,.38)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(95,99,104)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(32,33,36)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(23,78,166)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-t08AT-Bz112c{fill:rgba(95,99,104,.38)}.hqBSCb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-cTi5dd{color:rgb(95,99,104)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-cTi5dd{color:rgba(95,99,104,.38)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(197,34,31)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(165,14,14)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(197,34,31)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(197,34,31)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(165,14,14)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(197,34,31)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(165,14,14)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(217,48,37)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(165,14,14)}.hqBSCb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(217,48,37)}.hqBSCb .VfPpkd-TkwUic .VfPpkd-woaZLe::before,.hqBSCb .VfPpkd-TkwUic .VfPpkd-woaZLe::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.hqBSCb .VfPpkd-TkwUic:hover .VfPpkd-woaZLe::before,.hqBSCb .VfPpkd-TkwUic.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-woaZLe::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.hqBSCb .VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-woaZLe::before,.hqBSCb .VfPpkd-TkwUic:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-woaZLe::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.hqBSCb .VfPpkd-TkwUic:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-woaZLe::after{transition:opacity .15s linear}.hqBSCb .VfPpkd-TkwUic:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-woaZLe::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.hqBSCb .VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(128,134,139)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(32,33,36)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(26,115,232)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(60,64,67,.12)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(95,99,104)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(26,115,232)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(32,33,36)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(95,99,104,.38)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me)+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgb(95,99,104)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgba(95,99,104,.38)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(217,48,37)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover.VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(165,14,14)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-uusGie-fmcmS{color:rgb(60,64,67)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:rgba(60,64,67,.38)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(95,99,104)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(32,33,36)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(26,115,232)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-t08AT-Bz112c{fill:rgba(95,99,104,.38)}.ReCbLb:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-cTi5dd{color:rgb(95,99,104)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-cTi5dd{color:rgba(95,99,104,.38)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(217,48,37)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(165,14,14)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(217,48,37)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(217,48,37)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(165,14,14)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(217,48,37)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(165,14,14)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(197,34,31)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(165,14,14)}.ReCbLb.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(197,34,31)}.VfPpkd-BFbNVe-bF1uUb{position:absolute;border-radius:inherit;pointer-events:none;opacity:0;opacity:var(--mdc-elevation-overlay-opacity,0);transition:opacity .28s cubic-bezier(.4,0,.2,1);background-color:#fff;background-color:var(--mdc-elevation-overlay-color,#fff)}.VfPpkd-scr2fc{-moz-box-align:center;align-items:center;background:none;border:none;cursor:pointer;display:-moz-inline-box;display:inline-flex;flex-shrink:0;margin:0;outline:none;overflow:visible;padding:0;position:relative}.VfPpkd-scr2fc[hidden]{display:none}.VfPpkd-scr2fc:disabled{cursor:default;pointer-events:none}.VfPpkd-l6JLsf{overflow:hidden;position:relative;width:100%}.VfPpkd-l6JLsf::before,.VfPpkd-l6JLsf::after{border:1px solid transparent;border-radius:inherit;-moz-box-sizing:border-box;box-sizing:border-box;content:"";height:100%;left:0;position:absolute;width:100%}@media screen and (forced-colors:active){.VfPpkd-l6JLsf::before,.VfPpkd-l6JLsf::after{border-color:currentColor}}.VfPpkd-l6JLsf::before{transition:transform 75ms 0ms cubic-bezier(0,0,.2,1);transform:translateX(0)}.VfPpkd-l6JLsf::after{transition:transform 75ms 0ms cubic-bezier(.4,0,.6,1);transform:translateX(-100%)}[dir=rtl] .VfPpkd-l6JLsf::after,.VfPpkd-l6JLsf[dir=rtl]::after{transform:translateX(100%)}.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-l6JLsf::before{transition:transform 75ms 0ms cubic-bezier(.4,0,.6,1);transform:translateX(100%)}[dir=rtl] .VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-l6JLsf::before,.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-l6JLsf[dir=rtl]::before{transform:translateX(-100%)}.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-l6JLsf::after{transition:transform 75ms 0ms cubic-bezier(0,0,.2,1);transform:translateX(0)}.VfPpkd-uMhiad-u014N{height:100%;pointer-events:none;position:absolute;top:0;transition:transform 75ms 0ms cubic-bezier(.4,0,.2,1);left:0;right:auto;transform:translateX(0)}[dir=rtl] .VfPpkd-uMhiad-u014N,.VfPpkd-uMhiad-u014N[dir=rtl]{left:auto;right:0}.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-uMhiad-u014N{transform:translateX(100%)}[dir=rtl] .VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-uMhiad-u014N,.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-uMhiad-u014N[dir=rtl]{transform:translateX(-100%)}.VfPpkd-uMhiad{display:-moz-box;display:flex;pointer-events:auto;position:absolute;top:50%;transform:translateY(-50%);left:0;right:auto}[dir=rtl] .VfPpkd-uMhiad,.VfPpkd-uMhiad[dir=rtl]{left:auto;right:0}.VfPpkd-uMhiad::before,.VfPpkd-uMhiad::after{border:1px solid transparent;border-radius:inherit;-moz-box-sizing:border-box;box-sizing:border-box;content:"";width:100%;height:100%;left:0;position:absolute;top:0;transition:background-color 75ms 0ms cubic-bezier(.4,0,.2,1),border-color 75ms 0ms cubic-bezier(.4,0,.2,1);z-index:-1}@media screen and (forced-colors:active){.VfPpkd-uMhiad::before,.VfPpkd-uMhiad::after{border-color:currentColor}}.VfPpkd-VRSVNe{border-radius:inherit;bottom:0;left:0;position:absolute;right:0;top:0}.VfPpkd-BFbNVe-bF1uUb{bottom:0;left:0;right:0;top:0}.VfPpkd-Qsb3yd{left:50%;position:absolute;top:50%;transform:translate(-50%,-50%);z-index:-1}.VfPpkd-scr2fc:disabled .VfPpkd-Qsb3yd{display:none}.VfPpkd-lw9akd{height:100%;position:relative;width:100%;z-index:1}.VfPpkd-pafCAf{bottom:0;left:0;margin:auto;position:absolute;right:0;top:0;opacity:0;transition:opacity 30ms 0ms cubic-bezier(.4,0,1,1)}.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-pafCAf-OWXEXe-IT5dJd,.VfPpkd-scr2fc-OWXEXe-uqeOfd .VfPpkd-pafCAf-OWXEXe-Xhs9z{opacity:1;transition:opacity 45ms 30ms cubic-bezier(0,0,.2,1)}.VfPpkd-scr2fc{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-scr2fc .VfPpkd-Qsb3yd::before,.VfPpkd-scr2fc .VfPpkd-Qsb3yd::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-scr2fc .VfPpkd-Qsb3yd::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1}.VfPpkd-scr2fc .VfPpkd-Qsb3yd::after{z-index:0}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Qsb3yd::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Qsb3yd::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-Qsb3yd::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-Qsb3yd::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-Qsb3yd::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-scr2fc .VfPpkd-Qsb3yd::before,.VfPpkd-scr2fc .VfPpkd-Qsb3yd::after{top:0;left:0;width:100%;height:100%}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Qsb3yd::before,.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Qsb3yd::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0);width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Qsb3yd::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-scr2fc .VfPpkd-DVBDLb-LhBDec-sM5MNb{width:100%;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%)}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-DVBDLb-LhBDec,.VfPpkd-scr2fc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-DVBDLb-LhBDec{pointer-events:none;border:2px solid transparent;border-radius:6px;-moz-box-sizing:content-box;box-sizing:content-box;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-DVBDLb-LhBDec,.VfPpkd-scr2fc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-DVBDLb-LhBDec{border-color:CanvasText}}.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-DVBDLb-LhBDec::after,.VfPpkd-scr2fc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-DVBDLb-LhBDec::after{content:"";border:2px solid transparent;border-radius:8px;display:block;position:absolute;top:50%;left:50%;transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-scr2fc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-DVBDLb-LhBDec::after,.VfPpkd-scr2fc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-DVBDLb-LhBDec::after{border-color:CanvasText}}.LXctle{width:36px}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(26,115,232)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(23,78,166)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(23,78,166)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(23,78,166)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-uMhiad::after{background:rgb(60,64,67)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled .VfPpkd-uMhiad::after{background:rgb(95,99,104)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(32,33,36)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(32,33,36)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active .VfPpkd-uMhiad::after{background:rgb(32,33,36)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-uMhiad::after{background:rgb(60,64,67)}.LXctle .VfPpkd-uMhiad::before{background:rgb(255,255,255)}.LXctle:enabled .VfPpkd-VRSVNe{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15)}.LXctle:enabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.LXctle:enabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{background-color:transparent}.LXctle:disabled .VfPpkd-VRSVNe{box-shadow:none}.LXctle:disabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{opacity:0}.LXctle:disabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{background-color:transparent}.LXctle .VfPpkd-DVBDLb-LhBDec-sM5MNb,.LXctle .VfPpkd-uMhiad{height:20px}.LXctle:disabled .VfPpkd-uMhiad::after{opacity:.38}.LXctle .VfPpkd-uMhiad{border-radius:10px 10px 10px 10px}.LXctle .VfPpkd-uMhiad{width:20px}.LXctle .VfPpkd-uMhiad-u014N{width:calc(100% - 20px)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-pafCAf{fill:rgb(255,255,255)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-pafCAf{fill:rgb(255,255,255)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled .VfPpkd-pafCAf{fill:rgb(255,255,255)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-pafCAf{fill:rgb(255,255,255)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-lw9akd{opacity:.38}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-lw9akd{opacity:.38}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-pafCAf,.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd .VfPpkd-pafCAf{width:18px;height:18px}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(26,115,232)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(26,115,232)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(26,115,232)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(60,64,67)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(60,64,67)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(60,64,67)}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):hover .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe).VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Qsb3yd::before{opacity:.04}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Qsb3yd::before{transition-duration:75ms;opacity:.12}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Qsb3yd::after{transition:opacity .15s linear}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Qsb3yd::after{transition-duration:75ms;opacity:.1}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-switch-selected-pressed-state-layer-opacity,0.1)}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):hover .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe).VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Qsb3yd::before{opacity:.04}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Qsb3yd::before{transition-duration:75ms;opacity:.12}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Qsb3yd::after{transition:opacity .15s linear}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Qsb3yd::after{transition-duration:75ms;opacity:.1}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-switch-unselected-pressed-state-layer-opacity,0.1)}.LXctle .VfPpkd-Qsb3yd{height:48px;width:48px}.LXctle .VfPpkd-l6JLsf{height:14px}.LXctle:disabled .VfPpkd-l6JLsf{opacity:.12}.LXctle:enabled .VfPpkd-l6JLsf::after{background:rgb(138,180,248)}.LXctle:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:rgb(138,180,248)}.LXctle:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:rgb(138,180,248)}.LXctle:enabled:active .VfPpkd-l6JLsf::after{background:rgb(138,180,248)}.LXctle:disabled .VfPpkd-l6JLsf::after{background:rgb(60,64,67)}.LXctle:enabled .VfPpkd-l6JLsf::before{background:rgb(218,220,224)}.LXctle:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::before{background:rgb(218,220,224)}.LXctle:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::before{background:rgb(218,220,224)}.LXctle:enabled:active .VfPpkd-l6JLsf::before{background:rgb(218,220,224)}.LXctle:disabled .VfPpkd-l6JLsf::before{background:rgb(60,64,67)}.LXctle .VfPpkd-l6JLsf{border-radius:7px 7px 7px 7px}@media (-ms-high-contrast:active),screen and (forced-colors:active){.LXctle:disabled .VfPpkd-uMhiad::after{opacity:1}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-pafCAf{fill:ButtonText}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-pafCAf{fill:GrayText}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled .VfPpkd-pafCAf{fill:ButtonText}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-pafCAf{fill:GrayText}.LXctle.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-lw9akd{opacity:1}.LXctle.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-lw9akd{opacity:1}.LXctle:disabled .VfPpkd-l6JLsf{opacity:1}}.Ag4wUb.bFjUmb-Ysl7Fe,.Ag4wUb .bFjUmb-Ysl7Fe,.Ag4wUb.CNpREd.bFjUmb-Ysl7Fe,.Ag4wUb.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(232,240,254)}.Ag4wUb.bFjUmb-Wvd9Cc,.Ag4wUb .bFjUmb-Wvd9Cc,.Ag4wUb.CNpREd.bFjUmb-Wvd9Cc,.Ag4wUb.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(25,103,210)}.Ag4wUb.bFjUmb-Tvm9db,.Ag4wUb .bFjUmb-Tvm9db,.Ag4wUb.CNpREd.bFjUmb-Tvm9db,.Ag4wUb.CNpREd .bFjUmb-Tvm9db{background-color:rgb(23,78,166)}.Ag4wUb.yxp05b-Wvd9Cc,.Ag4wUb .yxp05b-Wvd9Cc,.Ag4wUb.CNpREd.yxp05b-Wvd9Cc,.Ag4wUb.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(25,103,210)}.Ag4wUb.VnOHwf-Ysl7Fe,.Ag4wUb .VnOHwf-Ysl7Fe,.Ag4wUb.CNpREd.VnOHwf-Ysl7Fe,.Ag4wUb.CNpREd .VnOHwf-Ysl7Fe{color:rgb(232,240,254);fill:rgb(232,240,254)}.Ag4wUb.VnOHwf-Wvd9Cc,.Ag4wUb .VnOHwf-Wvd9Cc,.Ag4wUb.CNpREd.VnOHwf-Wvd9Cc,.Ag4wUb.CNpREd .VnOHwf-Wvd9Cc{color:rgb(25,103,210);fill:rgb(25,103,210)}.Ag4wUb.VnOHwf-Tvm9db,.Ag4wUb .VnOHwf-Tvm9db,.Ag4wUb.CNpREd.VnOHwf-Tvm9db,.Ag4wUb.CNpREd .VnOHwf-Tvm9db{color:rgb(23,78,166);fill:rgb(23,78,166)}.Ag4wUb.eL9Cfb,.Ag4wUb .eL9Cfb,.Ag4wUb.L5mE7d,.Ag4wUb .L5mE7d,.Ag4wUb.eL9Cfb:hover,.Ag4wUb .eL9Cfb:hover,.Ag4wUb.eL9Cfb:focus,.Ag4wUb .eL9Cfb:focus,.Ag4wUb.CNpREd.eL9Cfb,.Ag4wUb.CNpREd .eL9Cfb,.Ag4wUb.CNpREd.L5mE7d,.Ag4wUb.CNpREd .L5mE7d,.Ag4wUb.CNpREd.eL9Cfb:hover,.Ag4wUb.CNpREd .eL9Cfb:hover,.Ag4wUb.CNpREd.eL9Cfb:focus,.Ag4wUb.CNpREd .eL9Cfb:focus{color:rgb(23,78,166)}.Ag4wUb.L5mE7d:hover,.Ag4wUb .L5mE7d:hover,.Ag4wUb.L5mE7d:focus,.Ag4wUb .L5mE7d:focus,.Ag4wUb.L5mE7d:visited,.Ag4wUb .L5mE7d:visited,.Ag4wUb.CNpREd.L5mE7d:hover,.Ag4wUb.CNpREd .L5mE7d:hover,.Ag4wUb.CNpREd.L5mE7d:focus,.Ag4wUb.CNpREd .L5mE7d:focus,.Ag4wUb.CNpREd.L5mE7d:visited,.Ag4wUb.CNpREd .L5mE7d:visited{color:rgb(25,103,210)}.Ag4wUb .VUoKZ{background-color:rgb(232,240,254)}.Ag4wUb .TRHLAc{background-color:rgb(25,103,210)}.Ag4wUb .tgNIJf-Ysl7Fe:focus{border-color:rgb(232,240,254)}.Ag4wUb .cjzpkc-Wvd9Cc:focus-within,.Ag4wUb .tgNIJf-Wvd9Cc:focus{border-color:rgb(25,103,210)}.Ag4wUb .u3bW4e .zZN2Lb-Wvd9Cc,.Ag4wUb .zZN2Lb-Wvd9Cc:focus,.Ag4wUb .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(25,103,210)}.Ag4wUb .P3W0Dd-Ysl7Fe:focus,.Ag4wUb.maXJsd:focus .P3W0Dd-Ysl7Fe,.Ag4wUb .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(232,240,254)}.Ag4wUb .VBEdtc-Wvd9Cc:hover,.Ag4wUb.MymH0d:hover .VBEdtc-Wvd9Cc,.Ag4wUb .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(25,103,210)}.Ag4wUb.MymH0d:hover .UISY8d-Tvm9db,.Ag4wUb.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.Ag4wUb .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(25,103,210)}.Ag4wUb .UISY8d-Ysl7Fe:hover,.Ag4wUb.MymH0d:hover .UISY8d-Ysl7Fe,.Ag4wUb .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(232,240,254)}.Ag4wUb .mxmXhf{color:rgb(23,78,166);fill:rgb(23,78,166)}.Ag4wUb .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.Ag4wUb .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.Ag4wUb .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.Ag4wUb .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.Ag4wUb .ZoT1D:focus-within.boxOzd,.Ag4wUb .ZoT1D:focus-within.idtp4e,.Ag4wUb .ZoT1D :focus-within.boxOzd,.Ag4wUb .ZoT1D :focus-within.idtp4e{background-color:rgb(232,240,254)}.Ag4wUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.Ag4wUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.Ag4wUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.Ag4wUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.Ag4wUb .ZoT1D:hover.j6KDAd,.Ag4wUb .ZoT1D:hover.idtp4e,.Ag4wUb .ZoT1D:hover .j6KDAd,.Ag4wUb .ZoT1D:hover .idtp4e{background-color:rgb(232,240,254)}.Ag4wUb .OGhwGf:hover,.Ag4wUb .OGhwGf:focus{color:rgb(23,78,166)}.Ag4wUb .ra2NV,.Ag4wUb.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(25,103,210),transparent)}.Ag4wUb .eumXzf:after{border-color:rgb(23,78,166)}.Ag4wUb .zKHdkd .cXrdqd,.Ag4wUb .kPBwDb{background-color:rgb(25,103,210)}.Ag4wUb .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.Ag4wUb .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(25,103,210)}.Ag4wUb .bkIpNd .uHMk6b{border-color:rgb(232,240,254)}.Ag4wUb .zJKIV .nQOrEb,.Ag4wUb .zJKIV.RDPZE .nQOrEb,.Ag4wUb .zJKIV.N2RpBe .Id5V1,.Ag4wUb .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(25,103,210)}.Ag4wUb .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(25,103,210);opacity:.5}.Ag4wUb .zJKIV.i9xfbb>.MbhUzd,.Ag4wUb .zJKIV.u3bW4e>.MbhUzd,.Ag4wUb .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.Ag4wUb .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(232,240,254)}.Ag4wUb .HQ8yf:not(.RDPZE),.Ag4wUb .HQ8yf:not(.RDPZE) a{color:rgb(25,103,210)}.Ag4wUb .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(25,103,210,.15)}.Ag4wUb .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(25,103,210,.25),rgba(25,103,210,.25) 80%,rgb(25,103,210) 100%)}.Ag4wUb .uO32ac,.Ag4wUb .ypv4re{border-bottom:1px solid rgb(25,103,210)}.Ag4wUb .DqwBN:not(.RDPZE) .TpQm9d,.Ag4wUb .l3F1ye:not(.RDPZE) .TpQm9d,.Ag4wUb .YhQJj:not(.RDPZE) .TpQm9d,.Ag4wUb .K2V86d:not(.RDPZE) .TpQm9d,.Ag4wUb .An19kf:not(.RDPZE) .TpQm9d{color:rgb(23,78,166);fill:rgb(23,78,166)}.Ag4wUb .DqwBN .TpQm9d,.Ag4wUb .YhQJj .TpQm9d,.Ag4wUb .K2V86d .TpQm9d,.Ag4wUb .l3F1ye .TpQm9d,.Ag4wUb .An19kf .TpQm9d{color:rgb(23,78,166);fill:rgb(23,78,166)}.Ag4wUb .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(138,180,248);fill:rgb(138,180,248)}.Ag4wUb .QkA63b:not(.RDPZE),.Ag4wUb .Y5sE8d:not(.RDPZE){background-color:rgb(23,78,166)}.Ag4wUb .An19kf:not(.RDPZE){background-color:rgb(232,240,254)}.Ag4wUb .QkA63b:not(.RDPZE):hover,.Ag4wUb .Y5sE8d:not(.RDPZE):hover,.Ag4wUb .QkA63b:not(.RDPZE).u3bW4e,.Ag4wUb .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(23,78,166,.2),0 1px 1px 0 rgba(23,78,166,.14),0 1px 3px 0 rgba(23,78,166,.12)}.Ag4wUb .QkA63b:not(.RDPZE).iWO5td,.Ag4wUb .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(23,78,166,.2),0 6px 10px 0 rgba(23,78,166,.14),0 1px 18px 0 rgba(23,78,166,.12)}.Ag4wUb .DqwBN:not(.RDPZE),.Ag4wUb .YhQJj:not(.RDPZE),.Ag4wUb .K2V86d:not(.RDPZE),.Ag4wUb .l3F1ye:not(.RDPZE),.Ag4wUb .An19kf:not(.RDPZE),.Ag4wUb .BEAGS:not(.RDPZE),.Ag4wUb .AeAAkf:not(.RDPZE){color:rgb(23,78,166)}.Ag4wUb .l3F1ye.j6PN2:not(.RDPZE){color:rgb(138,180,248)}.Ag4wUb .wwnMtb:not(.RDPZE),.Ag4wUb .OZ6W0d:not(.RDPZE){color:rgb(23,78,166);fill:rgb(23,78,166)}.Ag4wUb .wwnMtb:not(.RDPZE):hover,.Ag4wUb .OZ6W0d:not(.RDPZE):hover{background-color:rgba(23,78,166,.08)}.Ag4wUb .wwnMtb:not(.RDPZE).u3bW4e,.Ag4wUb .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(23,78,166,.12)}.Ag4wUb .wwnMtb:not(.RDPZE).u3bW4e:hover,.Ag4wUb .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(23,78,166,.16)}.Ag4wUb .BEAGS.iWO5td,.Ag4wUb .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(23,78,166,.2),0 1px 1px 0 rgba(23,78,166,.14),0 1px 3px 0 rgba(23,78,166,.12)}.Ag4wUb .DqwBN .MbhUzd,.Ag4wUb .YhQJj .MbhUzd,.Ag4wUb .K2V86d .MbhUzd,.Ag4wUb .l3F1ye .MbhUzd,.Ag4wUb .BEAGS .MbhUzd,.Ag4wUb .AeAAkf .MbhUzd,.Ag4wUb .An19kf .MbhUzd,.Ag4wUb .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(23,78,166,.16),rgba(23,78,166,.16) 80%,rgba(23,78,166,0) 100%)}.Ag4wUb .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(138,180,248,.16),rgba(138,180,248,.16) 80%,rgba(138,180,248,0) 100%)}.Ag4wUb .AeAAkf:not(.RDPZE) .CeoRYc,.Ag4wUb .BEAGS:not(.RDPZE) .CeoRYc,.Ag4wUb .An19kf:not(.RDPZE) .CeoRYc,.Ag4wUb .l3F1ye:not(.RDPZE) .CeoRYc,.Ag4wUb .YhQJj:not(.RDPZE) .CeoRYc,.Ag4wUb .K2V86d:not(.RDPZE) .CeoRYc,.Ag4wUb .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(23,78,166)}.Ag4wUb .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(138,180,248)}.Ag4wUb .AeAAkf:not(.RDPZE):hover,.Ag4wUb .AeAAkf:not(.RDPZE).u3bW4e,.Ag4wUb .BEAGS:not(.RDPZE):hover,.Ag4wUb .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(25,103,210,.2)}.Ag4wUb .DqwBN:not(.RDPZE):hover .CeoRYc,.Ag4wUb .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.Ag4wUb .YhQJj:not(.RDPZE):hover .CeoRYc,.Ag4wUb .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.Ag4wUb .K2V86d:not(.RDPZE):hover .CeoRYc,.Ag4wUb .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.Ag4wUb .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.Ag4wUb .l3F1ye:not(.RDPZE):hover .CeoRYc,.Ag4wUb .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(25,103,210)}.Ag4wUb .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.Ag4wUb .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(138,180,248)}.Ag4wUb .aiSeRd:not(.RDPZE).N2RpBe,.Ag4wUb .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(25,103,210)}.Ag4wUb .aiSeRd:not(.RDPZE):hover .MbhUzd,.Ag4wUb .aiSeRd:not(.RDPZE):focus .MbhUzd,.Ag4wUb .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.Ag4wUb .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(23,78,166,.08)}.Ag4wUb .d7L4fc:hover .hYsg7c,.Ag4wUb .NtlN8c:hover .hYsg7c{border-color:rgb(232,240,254)}.Ag4wUb .d7L4fc:hover .MbhUzd,.Ag4wUb .NtlN8c:hover .MbhUzd{background-color:rgba(23,78,166,.04)}.Ag4wUb .d7L4fc .hYsg7c .nQOrEb,.Ag4wUb .d7L4fc .hYsg7c.RDPZE .nQOrEb,.Ag4wUb .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(25,103,210)}.Ag4wUb .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.Ag4wUb .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(23,78,166,.08)}.Ag4wUb .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(25,103,210)}.Ag4wUb .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#5f9bec}.Ag4wUb .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(25,103,210,.3)}.Ag4wUb .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#bbd4f7}.Ag4wUb .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(25,103,210,.04)}.Ag4wUb .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.Ag4wUb .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.Ag4wUb .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(25,103,210,.12)}.Ag4wUb .HyS0Qd:not(.RDPZE) .zHQkBf,.Ag4wUb .fWf7qe:not(.RDPZE) .tL9Q4c,.Ag4wUb .D3oBEe:not(.RDPZE) .zHQkBf,.Ag4wUb .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(25,103,210)}.Ag4wUb .HyS0Qd:not(.RDPZE) .cXrdqd,.Ag4wUb .fWf7qe:not(.RDPZE) .cXrdqd,.Ag4wUb .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(25,103,210)}.Ag4wUb .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.Ag4wUb .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(25,103,210)}.Ag4wUb .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.Ag4wUb .HyS0Qd input:not([disabled]):focus~.snByac,.Ag4wUb .fWf7qe:not(.RDPZE).u3bW4e .snByac,.Ag4wUb .D3oBEe:not(.RDPZE).u3bW4e .snByac,.Ag4wUb .D3oBEe input:not([disabled]):focus~.snByac,.Ag4wUb .AkVYk:not(.RDPZE).u3bW4e .snByac,.Ag4wUb .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(23,78,166)}.Ag4wUb .ybOdnf:not(.RDPZE).iWO5td,.Ag4wUb .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.Ag4wUb .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(232,240,254)}.Ag4wUb .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(25,103,210);fill:rgb(25,103,210)}.Ag4wUb .mRipsb{background-color:rgb(25,103,210)}.Ag4wUb .bJuVn.KKjvXb{background-color:rgb(23,78,166)}.Ag4wUb .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(23,78,166),transparent)}.Ag4wUb .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(23,78,166),transparent)}.Ag4wUb .bJuVn.u3bW4e.KKjvXb.KKjvXb,.Ag4wUb .bJuVn.KKjvXb.KKjvXb:hover{background-color:#1955b4}.Ag4wUb .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.Ag4wUb .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#1955b4,transparent)}.Ag4wUb .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.Ag4wUb .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#1955b4,transparent)}.Ag4wUb .pAlOFe{color:rgb(23,78,166);fill:rgb(23,78,166)}.Ag4wUb .bDxw8b:not(:disabled){background-color:rgb(23,78,166)}.Ag4wUb .FL3Khc:not(:disabled){color:rgb(23,78,166)}.Ag4wUb .FL3Khc:not(:disabled):hover{color:rgb(23,78,166)}.Ag4wUb .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Ag4wUb .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(23,78,166)}.Ag4wUb .FL3Khc .VfPpkd-Jh9lGc::before,.Ag4wUb .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(23,78,166)}.Ag4wUb .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Ag4wUb .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(23,78,166)}.Ag4wUb .n42Gr:not(:disabled){color:rgb(23,78,166)}.Ag4wUb .n42Gr:not(:disabled):hover{color:rgb(23,78,166)}.Ag4wUb .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Ag4wUb .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(23,78,166)}.Ag4wUb .n42Gr .VfPpkd-Jh9lGc::before,.Ag4wUb .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(23,78,166)}.Ag4wUb .J5y29e:not(:disabled){color:rgb(23,78,166)}.Ag4wUb .J5y29e:not(:disabled):hover{color:rgb(23,78,166)}.Ag4wUb .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Ag4wUb .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(23,78,166)}.Ag4wUb .J5y29e .VfPpkd-Jh9lGc::before,.Ag4wUb .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(23,78,166)}.Ag4wUb .LgeCif{color:rgb(23,78,166)}.Ag4wUb .LgeCif:disabled{color:rgba(60,64,67,.38)}.Ag4wUb .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.Ag4wUb .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(23,78,166)}.Ag4wUb .wlZwYd:not(:disabled){background-color:rgb(232,240,254)}.Ag4wUb .wlZwYd:not(:disabled){color:rgb(23,78,166)}.Ag4wUb .wlZwYd:not(:disabled):hover{color:rgb(23,78,166)}.Ag4wUb .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Ag4wUb .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(23,78,166)}.Ag4wUb .wlZwYd .VfPpkd-Jh9lGc::before,.Ag4wUb .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(23,78,166)}.Ag4wUb .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.Ag4wUb .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-icon-color,rgb(25,103,210))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FF1967D200000000FF1967D2{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-icon-color,rgb(25,103,210))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FF1967D200000000FF1967D2{0%,80%{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-icon-color,rgb(25,103,210))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.Ag4wUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FF1967D200000000FF1967D2}.Ag4wUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FF1967D200000000FF1967D2}.Ag4wUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.Ag4wUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(23,78,166);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(23,78,166));background-color:rgb(23,78,166);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(23,78,166))}.Ag4wUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6}.Ag4wUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6}.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(23,78,166);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(23,78,166));background-color:rgb(23,78,166);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(23,78,166))}.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6}.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6}.Ag4wUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.Ag4wUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(23,78,166);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(23,78,166));background-color:rgb(23,78,166);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(23,78,166))}@keyframes mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(23,78,166);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(23,78,166));background-color:rgb(23,78,166);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(23,78,166))}}@keyframes mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6{0%,80%{border-color:rgb(23,78,166);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(23,78,166));background-color:rgb(23,78,166);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(23,78,166))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.Ag4wUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF174EA600000000FF174EA6}.Ag4wUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Ag4wUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF174EA600000000FF174EA6}.Ag4wUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.Ag4wUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(23,78,166);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(23,78,166))}.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.Ag4wUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(23,78,166);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(23,78,166))}.Ag4wUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.Ag4wUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.Ag4wUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.Ag4wUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.Ag4wUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.Ag4wUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(23,78,166)}.Ag4wUb .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob:hover .VfPpkd-eHTEvd::before,.Ag4wUb .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(23,78,166)}.Ag4wUb .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(25,103,210)}.Ag4wUb .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.Ag4wUb .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(23,78,166)}.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(25,103,210)}.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(23,78,166)}.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(23,78,166)}.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(23,78,166)}.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(23,78,166)}.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(23,78,166)}.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.Ag4wUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(23,78,166)}.Ag4wUb .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#9fc0fb}.Ag4wUb .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#9fc0fb}.Ag4wUb .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#9fc0fb}.Ag4wUb .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#9fc0fb}.Ag4wUb .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.Ag4wUb .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(23,78,166)}.Ag4wUb .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(23,78,166)}.Ag4wUb .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(23,78,166)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(25,103,210)}.Ag4wUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.Ag4wUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(25,103,210)}.Ag4wUb .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.Ag4wUb .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(25,103,210);background-color:var(--mdc-ripple-color,rgb(25,103,210))}.Ag4wUb .U5B3me:not(:disabled){color:rgb(138,180,248)}.Ag4wUb .U5B3me:not(:disabled):hover{color:rgb(138,180,248)}.Ag4wUb .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Ag4wUb .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(138,180,248)}.Ag4wUb .U5B3me .VfPpkd-Jh9lGc::before,.Ag4wUb .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(138,180,248)}.Ag4wUb .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(23,78,166)}.ee1HBc.bFjUmb-Ysl7Fe,.ee1HBc .bFjUmb-Ysl7Fe,.ee1HBc.CNpREd.bFjUmb-Ysl7Fe,.ee1HBc.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(232,240,254)}.ee1HBc.bFjUmb-Wvd9Cc,.ee1HBc .bFjUmb-Wvd9Cc,.ee1HBc.CNpREd.bFjUmb-Wvd9Cc,.ee1HBc.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(66,133,244)}.ee1HBc.bFjUmb-Tvm9db,.ee1HBc .bFjUmb-Tvm9db,.ee1HBc.CNpREd.bFjUmb-Tvm9db,.ee1HBc.CNpREd .bFjUmb-Tvm9db{background-color:rgb(25,103,210)}.ee1HBc.yxp05b-Wvd9Cc,.ee1HBc .yxp05b-Wvd9Cc,.ee1HBc.CNpREd.yxp05b-Wvd9Cc,.ee1HBc.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(66,133,244)}.ee1HBc.VnOHwf-Ysl7Fe,.ee1HBc .VnOHwf-Ysl7Fe,.ee1HBc.CNpREd.VnOHwf-Ysl7Fe,.ee1HBc.CNpREd .VnOHwf-Ysl7Fe{color:rgb(232,240,254);fill:rgb(232,240,254)}.ee1HBc.VnOHwf-Wvd9Cc,.ee1HBc .VnOHwf-Wvd9Cc,.ee1HBc.CNpREd.VnOHwf-Wvd9Cc,.ee1HBc.CNpREd .VnOHwf-Wvd9Cc{color:rgb(66,133,244);fill:rgb(66,133,244)}.ee1HBc.VnOHwf-Tvm9db,.ee1HBc .VnOHwf-Tvm9db,.ee1HBc.CNpREd.VnOHwf-Tvm9db,.ee1HBc.CNpREd .VnOHwf-Tvm9db{color:rgb(25,103,210);fill:rgb(25,103,210)}.ee1HBc.eL9Cfb,.ee1HBc .eL9Cfb,.ee1HBc.L5mE7d,.ee1HBc .L5mE7d,.ee1HBc.eL9Cfb:hover,.ee1HBc .eL9Cfb:hover,.ee1HBc.eL9Cfb:focus,.ee1HBc .eL9Cfb:focus,.ee1HBc.CNpREd.eL9Cfb,.ee1HBc.CNpREd .eL9Cfb,.ee1HBc.CNpREd.L5mE7d,.ee1HBc.CNpREd .L5mE7d,.ee1HBc.CNpREd.eL9Cfb:hover,.ee1HBc.CNpREd .eL9Cfb:hover,.ee1HBc.CNpREd.eL9Cfb:focus,.ee1HBc.CNpREd .eL9Cfb:focus{color:rgb(25,103,210)}.ee1HBc.L5mE7d:hover,.ee1HBc .L5mE7d:hover,.ee1HBc.L5mE7d:focus,.ee1HBc .L5mE7d:focus,.ee1HBc.L5mE7d:visited,.ee1HBc .L5mE7d:visited,.ee1HBc.CNpREd.L5mE7d:hover,.ee1HBc.CNpREd .L5mE7d:hover,.ee1HBc.CNpREd.L5mE7d:focus,.ee1HBc.CNpREd .L5mE7d:focus,.ee1HBc.CNpREd.L5mE7d:visited,.ee1HBc.CNpREd .L5mE7d:visited{color:rgb(66,133,244)}.ee1HBc .VUoKZ{background-color:rgb(232,240,254)}.ee1HBc .TRHLAc{background-color:rgb(66,133,244)}.ee1HBc .tgNIJf-Ysl7Fe:focus{border-color:rgb(232,240,254)}.ee1HBc .cjzpkc-Wvd9Cc:focus-within,.ee1HBc .tgNIJf-Wvd9Cc:focus{border-color:rgb(66,133,244)}.ee1HBc .u3bW4e .zZN2Lb-Wvd9Cc,.ee1HBc .zZN2Lb-Wvd9Cc:focus,.ee1HBc .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(66,133,244)}.ee1HBc .P3W0Dd-Ysl7Fe:focus,.ee1HBc.maXJsd:focus .P3W0Dd-Ysl7Fe,.ee1HBc .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(232,240,254)}.ee1HBc .VBEdtc-Wvd9Cc:hover,.ee1HBc.MymH0d:hover .VBEdtc-Wvd9Cc,.ee1HBc .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(66,133,244)}.ee1HBc.MymH0d:hover .UISY8d-Tvm9db,.ee1HBc.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.ee1HBc .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(66,133,244)}.ee1HBc .UISY8d-Ysl7Fe:hover,.ee1HBc.MymH0d:hover .UISY8d-Ysl7Fe,.ee1HBc .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(232,240,254)}.ee1HBc .mxmXhf{color:rgb(25,103,210);fill:rgb(25,103,210)}.ee1HBc .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.ee1HBc .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.ee1HBc .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.ee1HBc .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.ee1HBc .ZoT1D:focus-within.boxOzd,.ee1HBc .ZoT1D:focus-within.idtp4e,.ee1HBc .ZoT1D :focus-within.boxOzd,.ee1HBc .ZoT1D :focus-within.idtp4e{background-color:rgb(232,240,254)}.ee1HBc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.ee1HBc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.ee1HBc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.ee1HBc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.ee1HBc .ZoT1D:hover.j6KDAd,.ee1HBc .ZoT1D:hover.idtp4e,.ee1HBc .ZoT1D:hover .j6KDAd,.ee1HBc .ZoT1D:hover .idtp4e{background-color:rgb(232,240,254)}.ee1HBc .OGhwGf:hover,.ee1HBc .OGhwGf:focus{color:rgb(25,103,210)}.ee1HBc .ra2NV,.ee1HBc.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(66,133,244),transparent)}.ee1HBc .eumXzf:after{border-color:rgb(25,103,210)}.ee1HBc .zKHdkd .cXrdqd,.ee1HBc .kPBwDb{background-color:rgb(66,133,244)}.ee1HBc .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.ee1HBc .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(66,133,244)}.ee1HBc .bkIpNd .uHMk6b{border-color:rgb(232,240,254)}.ee1HBc .zJKIV .nQOrEb,.ee1HBc .zJKIV.RDPZE .nQOrEb,.ee1HBc .zJKIV.N2RpBe .Id5V1,.ee1HBc .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(66,133,244)}.ee1HBc .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(66,133,244);opacity:.5}.ee1HBc .zJKIV.i9xfbb>.MbhUzd,.ee1HBc .zJKIV.u3bW4e>.MbhUzd,.ee1HBc .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.ee1HBc .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(232,240,254)}.ee1HBc .HQ8yf:not(.RDPZE),.ee1HBc .HQ8yf:not(.RDPZE) a{color:rgb(66,133,244)}.ee1HBc .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(66,133,244,.15)}.ee1HBc .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(66,133,244,.25),rgba(66,133,244,.25) 80%,rgb(66,133,244) 100%)}.ee1HBc .uO32ac,.ee1HBc .ypv4re{border-bottom:1px solid rgb(66,133,244)}.ee1HBc .DqwBN:not(.RDPZE) .TpQm9d,.ee1HBc .l3F1ye:not(.RDPZE) .TpQm9d,.ee1HBc .YhQJj:not(.RDPZE) .TpQm9d,.ee1HBc .K2V86d:not(.RDPZE) .TpQm9d,.ee1HBc .An19kf:not(.RDPZE) .TpQm9d{color:rgb(25,103,210);fill:rgb(25,103,210)}.ee1HBc .DqwBN .TpQm9d,.ee1HBc .YhQJj .TpQm9d,.ee1HBc .K2V86d .TpQm9d,.ee1HBc .l3F1ye .TpQm9d,.ee1HBc .An19kf .TpQm9d{color:rgb(25,103,210);fill:rgb(25,103,210)}.ee1HBc .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(138,180,248);fill:rgb(138,180,248)}.ee1HBc .QkA63b:not(.RDPZE),.ee1HBc .Y5sE8d:not(.RDPZE){background-color:rgb(25,103,210)}.ee1HBc .An19kf:not(.RDPZE){background-color:rgb(232,240,254)}.ee1HBc .QkA63b:not(.RDPZE):hover,.ee1HBc .Y5sE8d:not(.RDPZE):hover,.ee1HBc .QkA63b:not(.RDPZE).u3bW4e,.ee1HBc .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(25,103,210,.2),0 1px 1px 0 rgba(25,103,210,.14),0 1px 3px 0 rgba(25,103,210,.12)}.ee1HBc .QkA63b:not(.RDPZE).iWO5td,.ee1HBc .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(25,103,210,.2),0 6px 10px 0 rgba(25,103,210,.14),0 1px 18px 0 rgba(25,103,210,.12)}.ee1HBc .DqwBN:not(.RDPZE),.ee1HBc .YhQJj:not(.RDPZE),.ee1HBc .K2V86d:not(.RDPZE),.ee1HBc .l3F1ye:not(.RDPZE),.ee1HBc .An19kf:not(.RDPZE),.ee1HBc .BEAGS:not(.RDPZE),.ee1HBc .AeAAkf:not(.RDPZE){color:rgb(25,103,210)}.ee1HBc .l3F1ye.j6PN2:not(.RDPZE){color:rgb(138,180,248)}.ee1HBc .wwnMtb:not(.RDPZE),.ee1HBc .OZ6W0d:not(.RDPZE){color:rgb(25,103,210);fill:rgb(25,103,210)}.ee1HBc .wwnMtb:not(.RDPZE):hover,.ee1HBc .OZ6W0d:not(.RDPZE):hover{background-color:rgba(25,103,210,.08)}.ee1HBc .wwnMtb:not(.RDPZE).u3bW4e,.ee1HBc .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(25,103,210,.12)}.ee1HBc .wwnMtb:not(.RDPZE).u3bW4e:hover,.ee1HBc .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(25,103,210,.16)}.ee1HBc .BEAGS.iWO5td,.ee1HBc .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(25,103,210,.2),0 1px 1px 0 rgba(25,103,210,.14),0 1px 3px 0 rgba(25,103,210,.12)}.ee1HBc .DqwBN .MbhUzd,.ee1HBc .YhQJj .MbhUzd,.ee1HBc .K2V86d .MbhUzd,.ee1HBc .l3F1ye .MbhUzd,.ee1HBc .BEAGS .MbhUzd,.ee1HBc .AeAAkf .MbhUzd,.ee1HBc .An19kf .MbhUzd,.ee1HBc .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(25,103,210,.16),rgba(25,103,210,.16) 80%,rgba(25,103,210,0) 100%)}.ee1HBc .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(138,180,248,.16),rgba(138,180,248,.16) 80%,rgba(138,180,248,0) 100%)}.ee1HBc .AeAAkf:not(.RDPZE) .CeoRYc,.ee1HBc .BEAGS:not(.RDPZE) .CeoRYc,.ee1HBc .An19kf:not(.RDPZE) .CeoRYc,.ee1HBc .l3F1ye:not(.RDPZE) .CeoRYc,.ee1HBc .YhQJj:not(.RDPZE) .CeoRYc,.ee1HBc .K2V86d:not(.RDPZE) .CeoRYc,.ee1HBc .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(25,103,210)}.ee1HBc .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(138,180,248)}.ee1HBc .AeAAkf:not(.RDPZE):hover,.ee1HBc .AeAAkf:not(.RDPZE).u3bW4e,.ee1HBc .BEAGS:not(.RDPZE):hover,.ee1HBc .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(66,133,244,.2)}.ee1HBc .DqwBN:not(.RDPZE):hover .CeoRYc,.ee1HBc .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.ee1HBc .YhQJj:not(.RDPZE):hover .CeoRYc,.ee1HBc .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.ee1HBc .K2V86d:not(.RDPZE):hover .CeoRYc,.ee1HBc .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.ee1HBc .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.ee1HBc .l3F1ye:not(.RDPZE):hover .CeoRYc,.ee1HBc .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(66,133,244)}.ee1HBc .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.ee1HBc .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(138,180,248)}.ee1HBc .aiSeRd:not(.RDPZE).N2RpBe,.ee1HBc .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(66,133,244)}.ee1HBc .aiSeRd:not(.RDPZE):hover .MbhUzd,.ee1HBc .aiSeRd:not(.RDPZE):focus .MbhUzd,.ee1HBc .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.ee1HBc .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(25,103,210,.08)}.ee1HBc .d7L4fc:hover .hYsg7c,.ee1HBc .NtlN8c:hover .hYsg7c{border-color:rgb(232,240,254)}.ee1HBc .d7L4fc:hover .MbhUzd,.ee1HBc .NtlN8c:hover .MbhUzd{background-color:rgba(25,103,210,.04)}.ee1HBc .d7L4fc .hYsg7c .nQOrEb,.ee1HBc .d7L4fc .hYsg7c.RDPZE .nQOrEb,.ee1HBc .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(66,133,244)}.ee1HBc .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.ee1HBc .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(25,103,210,.08)}.ee1HBc .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(66,133,244)}.ee1HBc .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#5692f5}.ee1HBc .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(66,133,244,.3)}.ee1HBc .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#b7d0fb}.ee1HBc .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(66,133,244,.04)}.ee1HBc .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.ee1HBc .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.ee1HBc .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(66,133,244,.12)}.ee1HBc .HyS0Qd:not(.RDPZE) .zHQkBf,.ee1HBc .fWf7qe:not(.RDPZE) .tL9Q4c,.ee1HBc .D3oBEe:not(.RDPZE) .zHQkBf,.ee1HBc .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(66,133,244)}.ee1HBc .HyS0Qd:not(.RDPZE) .cXrdqd,.ee1HBc .fWf7qe:not(.RDPZE) .cXrdqd,.ee1HBc .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(66,133,244)}.ee1HBc .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.ee1HBc .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(66,133,244)}.ee1HBc .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.ee1HBc .HyS0Qd input:not([disabled]):focus~.snByac,.ee1HBc .fWf7qe:not(.RDPZE).u3bW4e .snByac,.ee1HBc .D3oBEe:not(.RDPZE).u3bW4e .snByac,.ee1HBc .D3oBEe input:not([disabled]):focus~.snByac,.ee1HBc .AkVYk:not(.RDPZE).u3bW4e .snByac,.ee1HBc .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(25,103,210)}.ee1HBc .ybOdnf:not(.RDPZE).iWO5td,.ee1HBc .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.ee1HBc .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(232,240,254)}.ee1HBc .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(66,133,244);fill:rgb(66,133,244)}.ee1HBc .mRipsb{background-color:rgb(66,133,244)}.ee1HBc .bJuVn.KKjvXb{background-color:rgb(25,103,210)}.ee1HBc .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(25,103,210),transparent)}.ee1HBc .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(25,103,210),transparent)}.ee1HBc .bJuVn.u3bW4e.KKjvXb.KKjvXb,.ee1HBc .bJuVn.KKjvXb.KKjvXb:hover{background-color:#1a6dde}.ee1HBc .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.ee1HBc .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#1a6dde,transparent)}.ee1HBc .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.ee1HBc .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#1a6dde,transparent)}.ee1HBc .pAlOFe{color:rgb(25,103,210);fill:rgb(25,103,210)}.ee1HBc .bDxw8b:not(:disabled){background-color:rgb(25,103,210)}.ee1HBc .FL3Khc:not(:disabled){color:rgb(25,103,210)}.ee1HBc .FL3Khc:not(:disabled):hover{color:rgb(25,103,210)}.ee1HBc .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.ee1HBc .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(25,103,210)}.ee1HBc .FL3Khc .VfPpkd-Jh9lGc::before,.ee1HBc .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(25,103,210)}.ee1HBc .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.ee1HBc .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(25,103,210)}.ee1HBc .n42Gr:not(:disabled){color:rgb(25,103,210)}.ee1HBc .n42Gr:not(:disabled):hover{color:rgb(25,103,210)}.ee1HBc .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.ee1HBc .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(25,103,210)}.ee1HBc .n42Gr .VfPpkd-Jh9lGc::before,.ee1HBc .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(25,103,210)}.ee1HBc .J5y29e:not(:disabled){color:rgb(25,103,210)}.ee1HBc .J5y29e:not(:disabled):hover{color:rgb(25,103,210)}.ee1HBc .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.ee1HBc .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(25,103,210)}.ee1HBc .J5y29e .VfPpkd-Jh9lGc::before,.ee1HBc .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(25,103,210)}.ee1HBc .LgeCif{color:rgb(25,103,210)}.ee1HBc .LgeCif:disabled{color:rgba(60,64,67,.38)}.ee1HBc .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.ee1HBc .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(25,103,210)}.ee1HBc .wlZwYd:not(:disabled){background-color:rgb(232,240,254)}.ee1HBc .wlZwYd:not(:disabled){color:rgb(25,103,210)}.ee1HBc .wlZwYd:not(:disabled):hover{color:rgb(25,103,210)}.ee1HBc .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.ee1HBc .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(25,103,210)}.ee1HBc .wlZwYd .VfPpkd-Jh9lGc::before,.ee1HBc .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(25,103,210)}.ee1HBc .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.ee1HBc .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(66,133,244);border-color:var(--mdc-checkbox-selected-icon-color,rgb(66,133,244));background-color:rgb(66,133,244);background-color:var(--mdc-checkbox-selected-icon-color,rgb(66,133,244))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FF4285F400000000FF4285F4{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(66,133,244);border-color:var(--mdc-checkbox-selected-icon-color,rgb(66,133,244));background-color:rgb(66,133,244);background-color:var(--mdc-checkbox-selected-icon-color,rgb(66,133,244))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FF4285F400000000FF4285F4{0%,80%{border-color:rgb(66,133,244);border-color:var(--mdc-checkbox-selected-icon-color,rgb(66,133,244));background-color:rgb(66,133,244);background-color:var(--mdc-checkbox-selected-icon-color,rgb(66,133,244))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.ee1HBc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FF4285F400000000FF4285F4}.ee1HBc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FF4285F400000000FF4285F4}.ee1HBc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.ee1HBc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(25,103,210))}.ee1HBc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF1967D200000000FF1967D2}.ee1HBc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF1967D200000000FF1967D2}.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(25,103,210))}.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF1967D200000000FF1967D2}.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF1967D200000000FF1967D2}.ee1HBc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.ee1HBc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(25,103,210))}@keyframes mdc-checkbox-fade-in-background-FF202124FF1967D200000000FF1967D2{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(25,103,210))}}@keyframes mdc-checkbox-fade-out-background-FF202124FF1967D200000000FF1967D2{0%,80%{border-color:rgb(25,103,210);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(25,103,210));background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(25,103,210))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.ee1HBc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF1967D200000000FF1967D2}.ee1HBc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.ee1HBc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF1967D200000000FF1967D2}.ee1HBc .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.ee1HBc .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(25,103,210))}.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.ee1HBc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(25,103,210);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(25,103,210))}.ee1HBc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.ee1HBc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.ee1HBc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.ee1HBc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.ee1HBc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.ee1HBc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(25,103,210)}.ee1HBc .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob:hover .VfPpkd-eHTEvd::before,.ee1HBc .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(25,103,210)}.ee1HBc .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(66,133,244)}.ee1HBc .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.ee1HBc .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(25,103,210)}.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(66,133,244)}.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(25,103,210)}.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(25,103,210)}.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(25,103,210)}.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(25,103,210)}.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(25,103,210)}.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.ee1HBc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(25,103,210)}.ee1HBc .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#9fc0fb}.ee1HBc .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#9fc0fb}.ee1HBc .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#9fc0fb}.ee1HBc .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#9fc0fb}.ee1HBc .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.ee1HBc .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(25,103,210)}.ee1HBc .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(25,103,210)}.ee1HBc .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(25,103,210)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(66,133,244)}.ee1HBc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.ee1HBc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(66,133,244)}.ee1HBc .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.ee1HBc .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(66,133,244);background-color:var(--mdc-ripple-color,rgb(66,133,244))}.ee1HBc .U5B3me:not(:disabled){color:rgb(138,180,248)}.ee1HBc .U5B3me:not(:disabled):hover{color:rgb(138,180,248)}.ee1HBc .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.ee1HBc .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(138,180,248)}.ee1HBc .U5B3me .VfPpkd-Jh9lGc::before,.ee1HBc .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(138,180,248)}.ee1HBc .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(25,103,210)}.UvHKof.bFjUmb-Ysl7Fe,.UvHKof .bFjUmb-Ysl7Fe,.UvHKof.CNpREd.bFjUmb-Ysl7Fe,.UvHKof.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(241,243,244)}.UvHKof.bFjUmb-Wvd9Cc,.UvHKof .bFjUmb-Wvd9Cc,.UvHKof.CNpREd.bFjUmb-Wvd9Cc,.UvHKof.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(95,99,104)}.UvHKof.bFjUmb-Tvm9db,.UvHKof .bFjUmb-Tvm9db,.UvHKof.CNpREd.bFjUmb-Tvm9db,.UvHKof.CNpREd .bFjUmb-Tvm9db{background-color:rgb(32,33,36)}.UvHKof.yxp05b-Wvd9Cc,.UvHKof .yxp05b-Wvd9Cc,.UvHKof.CNpREd.yxp05b-Wvd9Cc,.UvHKof.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(95,99,104)}.UvHKof.VnOHwf-Ysl7Fe,.UvHKof .VnOHwf-Ysl7Fe,.UvHKof.CNpREd.VnOHwf-Ysl7Fe,.UvHKof.CNpREd .VnOHwf-Ysl7Fe{color:rgb(241,243,244);fill:rgb(241,243,244)}.UvHKof.VnOHwf-Wvd9Cc,.UvHKof .VnOHwf-Wvd9Cc,.UvHKof.CNpREd.VnOHwf-Wvd9Cc,.UvHKof.CNpREd .VnOHwf-Wvd9Cc{color:rgb(95,99,104);fill:rgb(95,99,104)}.UvHKof.VnOHwf-Tvm9db,.UvHKof .VnOHwf-Tvm9db,.UvHKof.CNpREd.VnOHwf-Tvm9db,.UvHKof.CNpREd .VnOHwf-Tvm9db{color:rgb(32,33,36);fill:rgb(32,33,36)}.UvHKof.eL9Cfb,.UvHKof .eL9Cfb,.UvHKof.L5mE7d,.UvHKof .L5mE7d,.UvHKof.eL9Cfb:hover,.UvHKof .eL9Cfb:hover,.UvHKof.eL9Cfb:focus,.UvHKof .eL9Cfb:focus,.UvHKof.CNpREd.eL9Cfb,.UvHKof.CNpREd .eL9Cfb,.UvHKof.CNpREd.L5mE7d,.UvHKof.CNpREd .L5mE7d,.UvHKof.CNpREd.eL9Cfb:hover,.UvHKof.CNpREd .eL9Cfb:hover,.UvHKof.CNpREd.eL9Cfb:focus,.UvHKof.CNpREd .eL9Cfb:focus{color:rgb(32,33,36)}.UvHKof.L5mE7d:hover,.UvHKof .L5mE7d:hover,.UvHKof.L5mE7d:focus,.UvHKof .L5mE7d:focus,.UvHKof.L5mE7d:visited,.UvHKof .L5mE7d:visited,.UvHKof.CNpREd.L5mE7d:hover,.UvHKof.CNpREd .L5mE7d:hover,.UvHKof.CNpREd.L5mE7d:focus,.UvHKof.CNpREd .L5mE7d:focus,.UvHKof.CNpREd.L5mE7d:visited,.UvHKof.CNpREd .L5mE7d:visited{color:rgb(95,99,104)}.UvHKof .VUoKZ{background-color:rgb(241,243,244)}.UvHKof .TRHLAc{background-color:rgb(95,99,104)}.UvHKof .tgNIJf-Ysl7Fe:focus{border-color:rgb(241,243,244)}.UvHKof .cjzpkc-Wvd9Cc:focus-within,.UvHKof .tgNIJf-Wvd9Cc:focus{border-color:rgb(95,99,104)}.UvHKof .u3bW4e .zZN2Lb-Wvd9Cc,.UvHKof .zZN2Lb-Wvd9Cc:focus,.UvHKof .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(95,99,104)}.UvHKof .P3W0Dd-Ysl7Fe:focus,.UvHKof.maXJsd:focus .P3W0Dd-Ysl7Fe,.UvHKof .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(241,243,244)}.UvHKof .VBEdtc-Wvd9Cc:hover,.UvHKof.MymH0d:hover .VBEdtc-Wvd9Cc,.UvHKof .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(95,99,104)}.UvHKof.MymH0d:hover .UISY8d-Tvm9db,.UvHKof.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.UvHKof .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(95,99,104)}.UvHKof .UISY8d-Ysl7Fe:hover,.UvHKof.MymH0d:hover .UISY8d-Ysl7Fe,.UvHKof .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(241,243,244)}.UvHKof .mxmXhf{color:rgb(32,33,36);fill:rgb(32,33,36)}.UvHKof .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.UvHKof .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.UvHKof .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.UvHKof .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.UvHKof .ZoT1D:focus-within.boxOzd,.UvHKof .ZoT1D:focus-within.idtp4e,.UvHKof .ZoT1D :focus-within.boxOzd,.UvHKof .ZoT1D :focus-within.idtp4e{background-color:rgb(241,243,244)}.UvHKof .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.UvHKof .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.UvHKof .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.UvHKof .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.UvHKof .ZoT1D:hover.j6KDAd,.UvHKof .ZoT1D:hover.idtp4e,.UvHKof .ZoT1D:hover .j6KDAd,.UvHKof .ZoT1D:hover .idtp4e{background-color:rgb(241,243,244)}.UvHKof .OGhwGf:hover,.UvHKof .OGhwGf:focus{color:rgb(32,33,36)}.UvHKof .ra2NV,.UvHKof.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(95,99,104),transparent)}.UvHKof .eumXzf:after{border-color:rgb(32,33,36)}.UvHKof .zKHdkd .cXrdqd,.UvHKof .kPBwDb{background-color:rgb(95,99,104)}.UvHKof .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.UvHKof .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(95,99,104)}.UvHKof .bkIpNd .uHMk6b{border-color:rgb(241,243,244)}.UvHKof .zJKIV .nQOrEb,.UvHKof .zJKIV.RDPZE .nQOrEb,.UvHKof .zJKIV.N2RpBe .Id5V1,.UvHKof .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(95,99,104)}.UvHKof .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(95,99,104);opacity:.5}.UvHKof .zJKIV.i9xfbb>.MbhUzd,.UvHKof .zJKIV.u3bW4e>.MbhUzd,.UvHKof .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.UvHKof .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(241,243,244)}.UvHKof .HQ8yf:not(.RDPZE),.UvHKof .HQ8yf:not(.RDPZE) a{color:rgb(95,99,104)}.UvHKof .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(95,99,104,.15)}.UvHKof .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(95,99,104,.25),rgba(95,99,104,.25) 80%,rgb(95,99,104) 100%)}.UvHKof .uO32ac,.UvHKof .ypv4re{border-bottom:1px solid rgb(95,99,104)}.UvHKof .DqwBN:not(.RDPZE) .TpQm9d,.UvHKof .l3F1ye:not(.RDPZE) .TpQm9d,.UvHKof .YhQJj:not(.RDPZE) .TpQm9d,.UvHKof .K2V86d:not(.RDPZE) .TpQm9d,.UvHKof .An19kf:not(.RDPZE) .TpQm9d{color:rgb(32,33,36);fill:rgb(32,33,36)}.UvHKof .DqwBN .TpQm9d,.UvHKof .YhQJj .TpQm9d,.UvHKof .K2V86d .TpQm9d,.UvHKof .l3F1ye .TpQm9d,.UvHKof .An19kf .TpQm9d{color:rgb(32,33,36);fill:rgb(32,33,36)}.UvHKof .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(218,220,224);fill:rgb(218,220,224)}.UvHKof .QkA63b:not(.RDPZE),.UvHKof .Y5sE8d:not(.RDPZE){background-color:rgb(32,33,36)}.UvHKof .An19kf:not(.RDPZE){background-color:rgb(241,243,244)}.UvHKof .QkA63b:not(.RDPZE):hover,.UvHKof .Y5sE8d:not(.RDPZE):hover,.UvHKof .QkA63b:not(.RDPZE).u3bW4e,.UvHKof .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(32,33,36,.2),0 1px 1px 0 rgba(32,33,36,.14),0 1px 3px 0 rgba(32,33,36,.12)}.UvHKof .QkA63b:not(.RDPZE).iWO5td,.UvHKof .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(32,33,36,.2),0 6px 10px 0 rgba(32,33,36,.14),0 1px 18px 0 rgba(32,33,36,.12)}.UvHKof .DqwBN:not(.RDPZE),.UvHKof .YhQJj:not(.RDPZE),.UvHKof .K2V86d:not(.RDPZE),.UvHKof .l3F1ye:not(.RDPZE),.UvHKof .An19kf:not(.RDPZE),.UvHKof .BEAGS:not(.RDPZE),.UvHKof .AeAAkf:not(.RDPZE){color:rgb(32,33,36)}.UvHKof .l3F1ye.j6PN2:not(.RDPZE){color:rgb(218,220,224)}.UvHKof .wwnMtb:not(.RDPZE),.UvHKof .OZ6W0d:not(.RDPZE){color:rgb(32,33,36);fill:rgb(32,33,36)}.UvHKof .wwnMtb:not(.RDPZE):hover,.UvHKof .OZ6W0d:not(.RDPZE):hover{background-color:rgba(32,33,36,.08)}.UvHKof .wwnMtb:not(.RDPZE).u3bW4e,.UvHKof .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(32,33,36,.12)}.UvHKof .wwnMtb:not(.RDPZE).u3bW4e:hover,.UvHKof .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(32,33,36,.16)}.UvHKof .BEAGS.iWO5td,.UvHKof .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(32,33,36,.2),0 1px 1px 0 rgba(32,33,36,.14),0 1px 3px 0 rgba(32,33,36,.12)}.UvHKof .DqwBN .MbhUzd,.UvHKof .YhQJj .MbhUzd,.UvHKof .K2V86d .MbhUzd,.UvHKof .l3F1ye .MbhUzd,.UvHKof .BEAGS .MbhUzd,.UvHKof .AeAAkf .MbhUzd,.UvHKof .An19kf .MbhUzd,.UvHKof .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(32,33,36,.16),rgba(32,33,36,.16) 80%,rgba(32,33,36,0) 100%)}.UvHKof .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(218,220,224,.16),rgba(218,220,224,.16) 80%,rgba(218,220,224,0) 100%)}.UvHKof .AeAAkf:not(.RDPZE) .CeoRYc,.UvHKof .BEAGS:not(.RDPZE) .CeoRYc,.UvHKof .An19kf:not(.RDPZE) .CeoRYc,.UvHKof .l3F1ye:not(.RDPZE) .CeoRYc,.UvHKof .YhQJj:not(.RDPZE) .CeoRYc,.UvHKof .K2V86d:not(.RDPZE) .CeoRYc,.UvHKof .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(32,33,36)}.UvHKof .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(218,220,224)}.UvHKof .AeAAkf:not(.RDPZE):hover,.UvHKof .AeAAkf:not(.RDPZE).u3bW4e,.UvHKof .BEAGS:not(.RDPZE):hover,.UvHKof .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(95,99,104,.2)}.UvHKof .DqwBN:not(.RDPZE):hover .CeoRYc,.UvHKof .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.UvHKof .YhQJj:not(.RDPZE):hover .CeoRYc,.UvHKof .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.UvHKof .K2V86d:not(.RDPZE):hover .CeoRYc,.UvHKof .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.UvHKof .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.UvHKof .l3F1ye:not(.RDPZE):hover .CeoRYc,.UvHKof .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(95,99,104)}.UvHKof .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.UvHKof .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(218,220,224)}.UvHKof .aiSeRd:not(.RDPZE).N2RpBe,.UvHKof .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(95,99,104)}.UvHKof .aiSeRd:not(.RDPZE):hover .MbhUzd,.UvHKof .aiSeRd:not(.RDPZE):focus .MbhUzd,.UvHKof .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.UvHKof .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(32,33,36,.08)}.UvHKof .d7L4fc:hover .hYsg7c,.UvHKof .NtlN8c:hover .hYsg7c{border-color:rgb(241,243,244)}.UvHKof .d7L4fc:hover .MbhUzd,.UvHKof .NtlN8c:hover .MbhUzd{background-color:rgba(32,33,36,.04)}.UvHKof .d7L4fc .hYsg7c .nQOrEb,.UvHKof .d7L4fc .hYsg7c.RDPZE .nQOrEb,.UvHKof .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(95,99,104)}.UvHKof .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.UvHKof .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(32,33,36,.08)}.UvHKof .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(95,99,104)}.UvHKof .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#a2a5aa}.UvHKof .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(95,99,104,.3)}.UvHKof .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#d7d9da}.UvHKof .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(95,99,104,.04)}.UvHKof .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.UvHKof .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.UvHKof .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(95,99,104,.12)}.UvHKof .HyS0Qd:not(.RDPZE) .zHQkBf,.UvHKof .fWf7qe:not(.RDPZE) .tL9Q4c,.UvHKof .D3oBEe:not(.RDPZE) .zHQkBf,.UvHKof .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(95,99,104)}.UvHKof .HyS0Qd:not(.RDPZE) .cXrdqd,.UvHKof .fWf7qe:not(.RDPZE) .cXrdqd,.UvHKof .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(95,99,104)}.UvHKof .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.UvHKof .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(95,99,104)}.UvHKof .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.UvHKof .HyS0Qd input:not([disabled]):focus~.snByac,.UvHKof .fWf7qe:not(.RDPZE).u3bW4e .snByac,.UvHKof .D3oBEe:not(.RDPZE).u3bW4e .snByac,.UvHKof .D3oBEe input:not([disabled]):focus~.snByac,.UvHKof .AkVYk:not(.RDPZE).u3bW4e .snByac,.UvHKof .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(32,33,36)}.UvHKof .ybOdnf:not(.RDPZE).iWO5td,.UvHKof .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.UvHKof .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(241,243,244)}.UvHKof .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(95,99,104);fill:rgb(95,99,104)}.UvHKof .mRipsb{background-color:rgb(95,99,104)}.UvHKof .bJuVn.KKjvXb{background-color:rgb(32,33,36)}.UvHKof .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(32,33,36),transparent)}.UvHKof .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(32,33,36),transparent)}.UvHKof .bJuVn.u3bW4e.KKjvXb.KKjvXb,.UvHKof .bJuVn.KKjvXb.KKjvXb:hover{background-color:#2a2c30}.UvHKof .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.UvHKof .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#2a2c30,transparent)}.UvHKof .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.UvHKof .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#2a2c30,transparent)}.UvHKof .pAlOFe{color:rgb(32,33,36);fill:rgb(32,33,36)}.UvHKof .bDxw8b:not(:disabled){background-color:rgb(32,33,36)}.UvHKof .FL3Khc:not(:disabled){color:rgb(32,33,36)}.UvHKof .FL3Khc:not(:disabled):hover{color:rgb(32,33,36)}.UvHKof .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.UvHKof .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36)}.UvHKof .FL3Khc .VfPpkd-Jh9lGc::before,.UvHKof .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36)}.UvHKof .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.UvHKof .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(32,33,36)}.UvHKof .n42Gr:not(:disabled){color:rgb(32,33,36)}.UvHKof .n42Gr:not(:disabled):hover{color:rgb(32,33,36)}.UvHKof .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.UvHKof .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36)}.UvHKof .n42Gr .VfPpkd-Jh9lGc::before,.UvHKof .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36)}.UvHKof .J5y29e:not(:disabled){color:rgb(32,33,36)}.UvHKof .J5y29e:not(:disabled):hover{color:rgb(32,33,36)}.UvHKof .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.UvHKof .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36)}.UvHKof .J5y29e .VfPpkd-Jh9lGc::before,.UvHKof .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36)}.UvHKof .LgeCif{color:rgb(32,33,36)}.UvHKof .LgeCif:disabled{color:rgba(60,64,67,.38)}.UvHKof .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.UvHKof .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(32,33,36)}.UvHKof .wlZwYd:not(:disabled){background-color:rgb(241,243,244)}.UvHKof .wlZwYd:not(:disabled){color:rgb(32,33,36)}.UvHKof .wlZwYd:not(:disabled):hover{color:rgb(32,33,36)}.UvHKof .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.UvHKof .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36)}.UvHKof .wlZwYd .VfPpkd-Jh9lGc::before,.UvHKof .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36)}.UvHKof .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.UvHKof .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.UvHKof .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.UvHKof .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-selected-icon-color,rgb(95,99,104));background-color:rgb(95,99,104);background-color:var(--mdc-checkbox-selected-icon-color,rgb(95,99,104))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FF5F636800000000FF5F6368{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-selected-icon-color,rgb(95,99,104));background-color:rgb(95,99,104);background-color:var(--mdc-checkbox-selected-icon-color,rgb(95,99,104))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FF5F636800000000FF5F6368{0%,80%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-selected-icon-color,rgb(95,99,104));background-color:rgb(95,99,104);background-color:var(--mdc-checkbox-selected-icon-color,rgb(95,99,104))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.UvHKof .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FF5F636800000000FF5F6368}.UvHKof .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FF5F636800000000FF5F6368}.UvHKof .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.UvHKof .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(32,33,36));background-color:rgb(32,33,36);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(32,33,36))}.UvHKof .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF20212400000000FF202124}.UvHKof .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF20212400000000FF202124}.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(32,33,36));background-color:rgb(32,33,36);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(32,33,36))}.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF20212400000000FF202124}.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF20212400000000FF202124}.UvHKof .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.UvHKof .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(32,33,36));background-color:rgb(32,33,36);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(32,33,36))}@keyframes mdc-checkbox-fade-in-background-FF202124FF20212400000000FF202124{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(32,33,36));background-color:rgb(32,33,36);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(32,33,36))}}@keyframes mdc-checkbox-fade-out-background-FF202124FF20212400000000FF202124{0%,80%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(32,33,36));background-color:rgb(32,33,36);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(32,33,36))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.UvHKof .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF20212400000000FF202124}.UvHKof .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.UvHKof .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF20212400000000FF202124}.UvHKof .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.UvHKof .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(32,33,36);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(32,33,36))}.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.UvHKof .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(32,33,36);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(32,33,36))}.UvHKof .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.UvHKof .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.UvHKof .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.UvHKof .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.UvHKof .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.UvHKof .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(32,33,36)}.UvHKof .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob:hover .VfPpkd-eHTEvd::before,.UvHKof .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(32,33,36)}.UvHKof .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(95,99,104)}.UvHKof .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.UvHKof .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(32,33,36)}.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(95,99,104)}.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(32,33,36)}.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(32,33,36)}.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(32,33,36)}.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(32,33,36)}.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(32,33,36)}.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.UvHKof .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(32,33,36)}.UvHKof .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#c6ced2}.UvHKof .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#c6ced2}.UvHKof .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#c6ced2}.UvHKof .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#c6ced2}.UvHKof .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(241,243,244)}.UvHKof .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(32,33,36)}.UvHKof .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(32,33,36)}.UvHKof .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(32,33,36)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(95,99,104)}.UvHKof .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.UvHKof .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(95,99,104)}.UvHKof .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.UvHKof .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(95,99,104);background-color:var(--mdc-ripple-color,rgb(95,99,104))}.UvHKof .U5B3me:not(:disabled){color:rgb(218,220,224)}.UvHKof .U5B3me:not(:disabled):hover{color:rgb(218,220,224)}.UvHKof .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.UvHKof .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(218,220,224)}.UvHKof .U5B3me .VfPpkd-Jh9lGc::before,.UvHKof .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(218,220,224)}.UvHKof .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(32,33,36)}.g2MItd.bFjUmb-Ysl7Fe,.g2MItd .bFjUmb-Ysl7Fe,.g2MItd.CNpREd.bFjUmb-Ysl7Fe,.g2MItd.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(254,239,227)}.g2MItd.bFjUmb-Wvd9Cc,.g2MItd .bFjUmb-Wvd9Cc,.g2MItd.CNpREd.bFjUmb-Wvd9Cc,.g2MItd.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(232,113,10)}.g2MItd.bFjUmb-Tvm9db,.g2MItd .bFjUmb-Tvm9db,.g2MItd.CNpREd.bFjUmb-Tvm9db,.g2MItd.CNpREd .bFjUmb-Tvm9db{background-color:rgb(194,100,1)}.g2MItd.yxp05b-Wvd9Cc,.g2MItd .yxp05b-Wvd9Cc,.g2MItd.CNpREd.yxp05b-Wvd9Cc,.g2MItd.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(232,113,10)}.g2MItd.VnOHwf-Ysl7Fe,.g2MItd .VnOHwf-Ysl7Fe,.g2MItd.CNpREd.VnOHwf-Ysl7Fe,.g2MItd.CNpREd .VnOHwf-Ysl7Fe{color:rgb(254,239,227);fill:rgb(254,239,227)}.g2MItd.VnOHwf-Wvd9Cc,.g2MItd .VnOHwf-Wvd9Cc,.g2MItd.CNpREd.VnOHwf-Wvd9Cc,.g2MItd.CNpREd .VnOHwf-Wvd9Cc{color:rgb(232,113,10);fill:rgb(232,113,10)}.g2MItd.VnOHwf-Tvm9db,.g2MItd .VnOHwf-Tvm9db,.g2MItd.CNpREd.VnOHwf-Tvm9db,.g2MItd.CNpREd .VnOHwf-Tvm9db{color:rgb(194,100,1);fill:rgb(194,100,1)}.g2MItd.eL9Cfb,.g2MItd .eL9Cfb,.g2MItd.L5mE7d,.g2MItd .L5mE7d,.g2MItd.eL9Cfb:hover,.g2MItd .eL9Cfb:hover,.g2MItd.eL9Cfb:focus,.g2MItd .eL9Cfb:focus,.g2MItd.CNpREd.eL9Cfb,.g2MItd.CNpREd .eL9Cfb,.g2MItd.CNpREd.L5mE7d,.g2MItd.CNpREd .L5mE7d,.g2MItd.CNpREd.eL9Cfb:hover,.g2MItd.CNpREd .eL9Cfb:hover,.g2MItd.CNpREd.eL9Cfb:focus,.g2MItd.CNpREd .eL9Cfb:focus{color:rgb(194,100,1)}.g2MItd.L5mE7d:hover,.g2MItd .L5mE7d:hover,.g2MItd.L5mE7d:focus,.g2MItd .L5mE7d:focus,.g2MItd.L5mE7d:visited,.g2MItd .L5mE7d:visited,.g2MItd.CNpREd.L5mE7d:hover,.g2MItd.CNpREd .L5mE7d:hover,.g2MItd.CNpREd.L5mE7d:focus,.g2MItd.CNpREd .L5mE7d:focus,.g2MItd.CNpREd.L5mE7d:visited,.g2MItd.CNpREd .L5mE7d:visited{color:rgb(232,113,10)}.g2MItd .VUoKZ{background-color:rgb(254,239,227)}.g2MItd .TRHLAc{background-color:rgb(232,113,10)}.g2MItd .tgNIJf-Ysl7Fe:focus{border-color:rgb(254,239,227)}.g2MItd .cjzpkc-Wvd9Cc:focus-within,.g2MItd .tgNIJf-Wvd9Cc:focus{border-color:rgb(232,113,10)}.g2MItd .u3bW4e .zZN2Lb-Wvd9Cc,.g2MItd .zZN2Lb-Wvd9Cc:focus,.g2MItd .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(232,113,10)}.g2MItd .P3W0Dd-Ysl7Fe:focus,.g2MItd.maXJsd:focus .P3W0Dd-Ysl7Fe,.g2MItd .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(254,239,227)}.g2MItd .VBEdtc-Wvd9Cc:hover,.g2MItd.MymH0d:hover .VBEdtc-Wvd9Cc,.g2MItd .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(232,113,10)}.g2MItd.MymH0d:hover .UISY8d-Tvm9db,.g2MItd.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.g2MItd .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(232,113,10)}.g2MItd .UISY8d-Ysl7Fe:hover,.g2MItd.MymH0d:hover .UISY8d-Ysl7Fe,.g2MItd .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(254,239,227)}.g2MItd .mxmXhf{color:rgb(194,100,1);fill:rgb(194,100,1)}.g2MItd .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.g2MItd .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.g2MItd .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.g2MItd .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.g2MItd .ZoT1D:focus-within.boxOzd,.g2MItd .ZoT1D:focus-within.idtp4e,.g2MItd .ZoT1D :focus-within.boxOzd,.g2MItd .ZoT1D :focus-within.idtp4e{background-color:rgb(254,239,227)}.g2MItd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.g2MItd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.g2MItd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.g2MItd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.g2MItd .ZoT1D:hover.j6KDAd,.g2MItd .ZoT1D:hover.idtp4e,.g2MItd .ZoT1D:hover .j6KDAd,.g2MItd .ZoT1D:hover .idtp4e{background-color:rgb(254,239,227)}.g2MItd .OGhwGf:hover,.g2MItd .OGhwGf:focus{color:rgb(194,100,1)}.g2MItd .ra2NV,.g2MItd.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(232,113,10),transparent)}.g2MItd .eumXzf:after{border-color:rgb(194,100,1)}.g2MItd .zKHdkd .cXrdqd,.g2MItd .kPBwDb{background-color:rgb(232,113,10)}.g2MItd .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.g2MItd .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(232,113,10)}.g2MItd .bkIpNd .uHMk6b{border-color:rgb(254,239,227)}.g2MItd .zJKIV .nQOrEb,.g2MItd .zJKIV.RDPZE .nQOrEb,.g2MItd .zJKIV.N2RpBe .Id5V1,.g2MItd .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(232,113,10)}.g2MItd .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(232,113,10);opacity:.5}.g2MItd .zJKIV.i9xfbb>.MbhUzd,.g2MItd .zJKIV.u3bW4e>.MbhUzd,.g2MItd .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.g2MItd .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(254,239,227)}.g2MItd .HQ8yf:not(.RDPZE),.g2MItd .HQ8yf:not(.RDPZE) a{color:rgb(232,113,10)}.g2MItd .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(232,113,10,.15)}.g2MItd .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(232,113,10,.25),rgba(232,113,10,.25) 80%,rgb(232,113,10) 100%)}.g2MItd .uO32ac,.g2MItd .ypv4re{border-bottom:1px solid rgb(232,113,10)}.g2MItd .DqwBN:not(.RDPZE) .TpQm9d,.g2MItd .l3F1ye:not(.RDPZE) .TpQm9d,.g2MItd .YhQJj:not(.RDPZE) .TpQm9d,.g2MItd .K2V86d:not(.RDPZE) .TpQm9d,.g2MItd .An19kf:not(.RDPZE) .TpQm9d{color:rgb(194,100,1);fill:rgb(194,100,1)}.g2MItd .DqwBN .TpQm9d,.g2MItd .YhQJj .TpQm9d,.g2MItd .K2V86d .TpQm9d,.g2MItd .l3F1ye .TpQm9d,.g2MItd .An19kf .TpQm9d{color:rgb(194,100,1);fill:rgb(194,100,1)}.g2MItd .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(252,173,112);fill:rgb(252,173,112)}.g2MItd .QkA63b:not(.RDPZE),.g2MItd .Y5sE8d:not(.RDPZE){background-color:rgb(194,100,1)}.g2MItd .An19kf:not(.RDPZE){background-color:rgb(254,239,227)}.g2MItd .QkA63b:not(.RDPZE):hover,.g2MItd .Y5sE8d:not(.RDPZE):hover,.g2MItd .QkA63b:not(.RDPZE).u3bW4e,.g2MItd .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(194,100,1,.2),0 1px 1px 0 rgba(194,100,1,.14),0 1px 3px 0 rgba(194,100,1,.12)}.g2MItd .QkA63b:not(.RDPZE).iWO5td,.g2MItd .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(194,100,1,.2),0 6px 10px 0 rgba(194,100,1,.14),0 1px 18px 0 rgba(194,100,1,.12)}.g2MItd .DqwBN:not(.RDPZE),.g2MItd .YhQJj:not(.RDPZE),.g2MItd .K2V86d:not(.RDPZE),.g2MItd .l3F1ye:not(.RDPZE),.g2MItd .An19kf:not(.RDPZE),.g2MItd .BEAGS:not(.RDPZE),.g2MItd .AeAAkf:not(.RDPZE){color:rgb(194,100,1)}.g2MItd .l3F1ye.j6PN2:not(.RDPZE){color:rgb(252,173,112)}.g2MItd .wwnMtb:not(.RDPZE),.g2MItd .OZ6W0d:not(.RDPZE){color:rgb(194,100,1);fill:rgb(194,100,1)}.g2MItd .wwnMtb:not(.RDPZE):hover,.g2MItd .OZ6W0d:not(.RDPZE):hover{background-color:rgba(194,100,1,.08)}.g2MItd .wwnMtb:not(.RDPZE).u3bW4e,.g2MItd .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(194,100,1,.12)}.g2MItd .wwnMtb:not(.RDPZE).u3bW4e:hover,.g2MItd .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(194,100,1,.16)}.g2MItd .BEAGS.iWO5td,.g2MItd .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(194,100,1,.2),0 1px 1px 0 rgba(194,100,1,.14),0 1px 3px 0 rgba(194,100,1,.12)}.g2MItd .DqwBN .MbhUzd,.g2MItd .YhQJj .MbhUzd,.g2MItd .K2V86d .MbhUzd,.g2MItd .l3F1ye .MbhUzd,.g2MItd .BEAGS .MbhUzd,.g2MItd .AeAAkf .MbhUzd,.g2MItd .An19kf .MbhUzd,.g2MItd .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(194,100,1,.16),rgba(194,100,1,.16) 80%,rgba(194,100,1,0) 100%)}.g2MItd .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(252,173,112,.16),rgba(252,173,112,.16) 80%,rgba(252,173,112,0) 100%)}.g2MItd .AeAAkf:not(.RDPZE) .CeoRYc,.g2MItd .BEAGS:not(.RDPZE) .CeoRYc,.g2MItd .An19kf:not(.RDPZE) .CeoRYc,.g2MItd .l3F1ye:not(.RDPZE) .CeoRYc,.g2MItd .YhQJj:not(.RDPZE) .CeoRYc,.g2MItd .K2V86d:not(.RDPZE) .CeoRYc,.g2MItd .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(194,100,1)}.g2MItd .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(252,173,112)}.g2MItd .AeAAkf:not(.RDPZE):hover,.g2MItd .AeAAkf:not(.RDPZE).u3bW4e,.g2MItd .BEAGS:not(.RDPZE):hover,.g2MItd .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(232,113,10,.2)}.g2MItd .DqwBN:not(.RDPZE):hover .CeoRYc,.g2MItd .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.g2MItd .YhQJj:not(.RDPZE):hover .CeoRYc,.g2MItd .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.g2MItd .K2V86d:not(.RDPZE):hover .CeoRYc,.g2MItd .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.g2MItd .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.g2MItd .l3F1ye:not(.RDPZE):hover .CeoRYc,.g2MItd .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(232,113,10)}.g2MItd .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.g2MItd .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(252,173,112)}.g2MItd .aiSeRd:not(.RDPZE).N2RpBe,.g2MItd .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(232,113,10)}.g2MItd .aiSeRd:not(.RDPZE):hover .MbhUzd,.g2MItd .aiSeRd:not(.RDPZE):focus .MbhUzd,.g2MItd .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.g2MItd .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(194,100,1,.08)}.g2MItd .d7L4fc:hover .hYsg7c,.g2MItd .NtlN8c:hover .hYsg7c{border-color:rgb(254,239,227)}.g2MItd .d7L4fc:hover .MbhUzd,.g2MItd .NtlN8c:hover .MbhUzd{background-color:rgba(194,100,1,.04)}.g2MItd .d7L4fc .hYsg7c .nQOrEb,.g2MItd .d7L4fc .hYsg7c.RDPZE .nQOrEb,.g2MItd .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(232,113,10)}.g2MItd .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.g2MItd .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(194,100,1,.08)}.g2MItd .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(232,113,10)}.g2MItd .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#f8a054}.g2MItd .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(232,113,10,.3)}.g2MItd .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#fcd6b6}.g2MItd .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(232,113,10,.04)}.g2MItd .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.g2MItd .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.g2MItd .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(232,113,10,.12)}.g2MItd .HyS0Qd:not(.RDPZE) .zHQkBf,.g2MItd .fWf7qe:not(.RDPZE) .tL9Q4c,.g2MItd .D3oBEe:not(.RDPZE) .zHQkBf,.g2MItd .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(232,113,10)}.g2MItd .HyS0Qd:not(.RDPZE) .cXrdqd,.g2MItd .fWf7qe:not(.RDPZE) .cXrdqd,.g2MItd .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(232,113,10)}.g2MItd .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.g2MItd .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(232,113,10)}.g2MItd .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.g2MItd .HyS0Qd input:not([disabled]):focus~.snByac,.g2MItd .fWf7qe:not(.RDPZE).u3bW4e .snByac,.g2MItd .D3oBEe:not(.RDPZE).u3bW4e .snByac,.g2MItd .D3oBEe input:not([disabled]):focus~.snByac,.g2MItd .AkVYk:not(.RDPZE).u3bW4e .snByac,.g2MItd .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(194,100,1)}.g2MItd .ybOdnf:not(.RDPZE).iWO5td,.g2MItd .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.g2MItd .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(254,239,227)}.g2MItd .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(232,113,10);fill:rgb(232,113,10)}.g2MItd .mRipsb{background-color:rgb(232,113,10)}.g2MItd .bJuVn.KKjvXb{background-color:rgb(194,100,1)}.g2MItd .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(194,100,1),transparent)}.g2MItd .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(194,100,1),transparent)}.g2MItd .bJuVn.u3bW4e.KKjvXb.KKjvXb,.g2MItd .bJuVn.KKjvXb.KKjvXb:hover{background-color:#d26c01}.g2MItd .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.g2MItd .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#d26c01,transparent)}.g2MItd .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.g2MItd .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#d26c01,transparent)}.g2MItd .pAlOFe{color:rgb(194,100,1);fill:rgb(194,100,1)}.g2MItd .bDxw8b:not(:disabled){background-color:rgb(194,100,1)}.g2MItd .FL3Khc:not(:disabled){color:rgb(194,100,1)}.g2MItd .FL3Khc:not(:disabled):hover{color:rgb(194,100,1)}.g2MItd .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.g2MItd .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(194,100,1)}.g2MItd .FL3Khc .VfPpkd-Jh9lGc::before,.g2MItd .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(194,100,1)}.g2MItd .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.g2MItd .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(194,100,1)}.g2MItd .n42Gr:not(:disabled){color:rgb(194,100,1)}.g2MItd .n42Gr:not(:disabled):hover{color:rgb(194,100,1)}.g2MItd .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.g2MItd .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(194,100,1)}.g2MItd .n42Gr .VfPpkd-Jh9lGc::before,.g2MItd .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(194,100,1)}.g2MItd .J5y29e:not(:disabled){color:rgb(194,100,1)}.g2MItd .J5y29e:not(:disabled):hover{color:rgb(194,100,1)}.g2MItd .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.g2MItd .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(194,100,1)}.g2MItd .J5y29e .VfPpkd-Jh9lGc::before,.g2MItd .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(194,100,1)}.g2MItd .LgeCif{color:rgb(194,100,1)}.g2MItd .LgeCif:disabled{color:rgba(60,64,67,.38)}.g2MItd .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.g2MItd .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(194,100,1)}.g2MItd .wlZwYd:not(:disabled){background-color:rgb(254,239,227)}.g2MItd .wlZwYd:not(:disabled){color:rgb(194,100,1)}.g2MItd .wlZwYd:not(:disabled):hover{color:rgb(194,100,1)}.g2MItd .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.g2MItd .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(194,100,1)}.g2MItd .wlZwYd .VfPpkd-Jh9lGc::before,.g2MItd .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(194,100,1)}.g2MItd .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.g2MItd .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.g2MItd .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.g2MItd .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(232,113,10);border-color:var(--mdc-checkbox-selected-icon-color,rgb(232,113,10));background-color:rgb(232,113,10);background-color:var(--mdc-checkbox-selected-icon-color,rgb(232,113,10))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FFE8710A00000000FFE8710A{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(232,113,10);border-color:var(--mdc-checkbox-selected-icon-color,rgb(232,113,10));background-color:rgb(232,113,10);background-color:var(--mdc-checkbox-selected-icon-color,rgb(232,113,10))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FFE8710A00000000FFE8710A{0%,80%{border-color:rgb(232,113,10);border-color:var(--mdc-checkbox-selected-icon-color,rgb(232,113,10));background-color:rgb(232,113,10);background-color:var(--mdc-checkbox-selected-icon-color,rgb(232,113,10))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.g2MItd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FFE8710A00000000FFE8710A}.g2MItd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FFE8710A00000000FFE8710A}.g2MItd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.g2MItd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(194,100,1);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(194,100,1));background-color:rgb(194,100,1);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(194,100,1))}.g2MItd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FFC2640100000000FFC26401}.g2MItd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FFC2640100000000FFC26401}.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(194,100,1);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(194,100,1));background-color:rgb(194,100,1);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(194,100,1))}.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FFC2640100000000FFC26401}.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FFC2640100000000FFC26401}.g2MItd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.g2MItd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(194,100,1);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(194,100,1));background-color:rgb(194,100,1);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(194,100,1))}@keyframes mdc-checkbox-fade-in-background-FF202124FFC2640100000000FFC26401{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(194,100,1);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(194,100,1));background-color:rgb(194,100,1);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(194,100,1))}}@keyframes mdc-checkbox-fade-out-background-FF202124FFC2640100000000FFC26401{0%,80%{border-color:rgb(194,100,1);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(194,100,1));background-color:rgb(194,100,1);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(194,100,1))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.g2MItd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FFC2640100000000FFC26401}.g2MItd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.g2MItd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FFC2640100000000FFC26401}.g2MItd .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.g2MItd .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(194,100,1);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(194,100,1))}.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.g2MItd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(194,100,1);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(194,100,1))}.g2MItd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.g2MItd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.g2MItd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.g2MItd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.g2MItd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.g2MItd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(194,100,1)}.g2MItd .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob:hover .VfPpkd-eHTEvd::before,.g2MItd .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(194,100,1)}.g2MItd .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(232,113,10)}.g2MItd .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.g2MItd .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(194,100,1)}.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(232,113,10)}.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(194,100,1)}.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(194,100,1)}.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(194,100,1)}.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(194,100,1)}.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(194,100,1)}.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.g2MItd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(194,100,1)}.g2MItd .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#fbc599}.g2MItd .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#fbc599}.g2MItd .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#fbc599}.g2MItd .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#fbc599}.g2MItd .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(254,239,227)}.g2MItd .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(194,100,1)}.g2MItd .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(194,100,1)}.g2MItd .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(194,100,1)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(232,113,10)}.g2MItd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.g2MItd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(232,113,10)}.g2MItd .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.g2MItd .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(232,113,10);background-color:var(--mdc-ripple-color,rgb(232,113,10))}.g2MItd .U5B3me:not(:disabled){color:rgb(252,173,112)}.g2MItd .U5B3me:not(:disabled):hover{color:rgb(252,173,112)}.g2MItd .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.g2MItd .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(252,173,112)}.g2MItd .U5B3me .VfPpkd-Jh9lGc::before,.g2MItd .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(252,173,112)}.g2MItd .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(194,100,1)}.S3aLQd.bFjUmb-Ysl7Fe,.S3aLQd .bFjUmb-Ysl7Fe,.S3aLQd.CNpREd.bFjUmb-Ysl7Fe,.S3aLQd.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(228,247,251)}.S3aLQd.bFjUmb-Wvd9Cc,.S3aLQd .bFjUmb-Wvd9Cc,.S3aLQd.CNpREd.bFjUmb-Wvd9Cc,.S3aLQd.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(18,158,175)}.S3aLQd.bFjUmb-Tvm9db,.S3aLQd .bFjUmb-Tvm9db,.S3aLQd.CNpREd.bFjUmb-Tvm9db,.S3aLQd.CNpREd .bFjUmb-Tvm9db{background-color:rgb(0,123,131)}.S3aLQd.yxp05b-Wvd9Cc,.S3aLQd .yxp05b-Wvd9Cc,.S3aLQd.CNpREd.yxp05b-Wvd9Cc,.S3aLQd.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(18,158,175)}.S3aLQd.VnOHwf-Ysl7Fe,.S3aLQd .VnOHwf-Ysl7Fe,.S3aLQd.CNpREd.VnOHwf-Ysl7Fe,.S3aLQd.CNpREd .VnOHwf-Ysl7Fe{color:rgb(228,247,251);fill:rgb(228,247,251)}.S3aLQd.VnOHwf-Wvd9Cc,.S3aLQd .VnOHwf-Wvd9Cc,.S3aLQd.CNpREd.VnOHwf-Wvd9Cc,.S3aLQd.CNpREd .VnOHwf-Wvd9Cc{color:rgb(18,158,175);fill:rgb(18,158,175)}.S3aLQd.VnOHwf-Tvm9db,.S3aLQd .VnOHwf-Tvm9db,.S3aLQd.CNpREd.VnOHwf-Tvm9db,.S3aLQd.CNpREd .VnOHwf-Tvm9db{color:rgb(0,123,131);fill:rgb(0,123,131)}.S3aLQd.eL9Cfb,.S3aLQd .eL9Cfb,.S3aLQd.L5mE7d,.S3aLQd .L5mE7d,.S3aLQd.eL9Cfb:hover,.S3aLQd .eL9Cfb:hover,.S3aLQd.eL9Cfb:focus,.S3aLQd .eL9Cfb:focus,.S3aLQd.CNpREd.eL9Cfb,.S3aLQd.CNpREd .eL9Cfb,.S3aLQd.CNpREd.L5mE7d,.S3aLQd.CNpREd .L5mE7d,.S3aLQd.CNpREd.eL9Cfb:hover,.S3aLQd.CNpREd .eL9Cfb:hover,.S3aLQd.CNpREd.eL9Cfb:focus,.S3aLQd.CNpREd .eL9Cfb:focus{color:rgb(0,123,131)}.S3aLQd.L5mE7d:hover,.S3aLQd .L5mE7d:hover,.S3aLQd.L5mE7d:focus,.S3aLQd .L5mE7d:focus,.S3aLQd.L5mE7d:visited,.S3aLQd .L5mE7d:visited,.S3aLQd.CNpREd.L5mE7d:hover,.S3aLQd.CNpREd .L5mE7d:hover,.S3aLQd.CNpREd.L5mE7d:focus,.S3aLQd.CNpREd .L5mE7d:focus,.S3aLQd.CNpREd.L5mE7d:visited,.S3aLQd.CNpREd .L5mE7d:visited{color:rgb(18,158,175)}.S3aLQd .VUoKZ{background-color:rgb(228,247,251)}.S3aLQd .TRHLAc{background-color:rgb(18,158,175)}.S3aLQd .tgNIJf-Ysl7Fe:focus{border-color:rgb(228,247,251)}.S3aLQd .cjzpkc-Wvd9Cc:focus-within,.S3aLQd .tgNIJf-Wvd9Cc:focus{border-color:rgb(18,158,175)}.S3aLQd .u3bW4e .zZN2Lb-Wvd9Cc,.S3aLQd .zZN2Lb-Wvd9Cc:focus,.S3aLQd .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(18,158,175)}.S3aLQd .P3W0Dd-Ysl7Fe:focus,.S3aLQd.maXJsd:focus .P3W0Dd-Ysl7Fe,.S3aLQd .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(228,247,251)}.S3aLQd .VBEdtc-Wvd9Cc:hover,.S3aLQd.MymH0d:hover .VBEdtc-Wvd9Cc,.S3aLQd .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(18,158,175)}.S3aLQd.MymH0d:hover .UISY8d-Tvm9db,.S3aLQd.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.S3aLQd .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(18,158,175)}.S3aLQd .UISY8d-Ysl7Fe:hover,.S3aLQd.MymH0d:hover .UISY8d-Ysl7Fe,.S3aLQd .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(228,247,251)}.S3aLQd .mxmXhf{color:rgb(0,123,131);fill:rgb(0,123,131)}.S3aLQd .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.S3aLQd .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.S3aLQd .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.S3aLQd .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.S3aLQd .ZoT1D:focus-within.boxOzd,.S3aLQd .ZoT1D:focus-within.idtp4e,.S3aLQd .ZoT1D :focus-within.boxOzd,.S3aLQd .ZoT1D :focus-within.idtp4e{background-color:rgb(228,247,251)}.S3aLQd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.S3aLQd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.S3aLQd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.S3aLQd .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.S3aLQd .ZoT1D:hover.j6KDAd,.S3aLQd .ZoT1D:hover.idtp4e,.S3aLQd .ZoT1D:hover .j6KDAd,.S3aLQd .ZoT1D:hover .idtp4e{background-color:rgb(228,247,251)}.S3aLQd .OGhwGf:hover,.S3aLQd .OGhwGf:focus{color:rgb(0,123,131)}.S3aLQd .ra2NV,.S3aLQd.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(18,158,175),transparent)}.S3aLQd .eumXzf:after{border-color:rgb(0,123,131)}.S3aLQd .zKHdkd .cXrdqd,.S3aLQd .kPBwDb{background-color:rgb(18,158,175)}.S3aLQd .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.S3aLQd .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(18,158,175)}.S3aLQd .bkIpNd .uHMk6b{border-color:rgb(228,247,251)}.S3aLQd .zJKIV .nQOrEb,.S3aLQd .zJKIV.RDPZE .nQOrEb,.S3aLQd .zJKIV.N2RpBe .Id5V1,.S3aLQd .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(18,158,175)}.S3aLQd .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(18,158,175);opacity:.5}.S3aLQd .zJKIV.i9xfbb>.MbhUzd,.S3aLQd .zJKIV.u3bW4e>.MbhUzd,.S3aLQd .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.S3aLQd .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(228,247,251)}.S3aLQd .HQ8yf:not(.RDPZE),.S3aLQd .HQ8yf:not(.RDPZE) a{color:rgb(18,158,175)}.S3aLQd .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(18,158,175,.15)}.S3aLQd .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(18,158,175,.25),rgba(18,158,175,.25) 80%,rgb(18,158,175) 100%)}.S3aLQd .uO32ac,.S3aLQd .ypv4re{border-bottom:1px solid rgb(18,158,175)}.S3aLQd .DqwBN:not(.RDPZE) .TpQm9d,.S3aLQd .l3F1ye:not(.RDPZE) .TpQm9d,.S3aLQd .YhQJj:not(.RDPZE) .TpQm9d,.S3aLQd .K2V86d:not(.RDPZE) .TpQm9d,.S3aLQd .An19kf:not(.RDPZE) .TpQm9d{color:rgb(0,123,131);fill:rgb(0,123,131)}.S3aLQd .DqwBN .TpQm9d,.S3aLQd .YhQJj .TpQm9d,.S3aLQd .K2V86d .TpQm9d,.S3aLQd .l3F1ye .TpQm9d,.S3aLQd .An19kf .TpQm9d{color:rgb(0,123,131);fill:rgb(0,123,131)}.S3aLQd .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(120,217,236);fill:rgb(120,217,236)}.S3aLQd .QkA63b:not(.RDPZE),.S3aLQd .Y5sE8d:not(.RDPZE){background-color:rgb(0,123,131)}.S3aLQd .An19kf:not(.RDPZE){background-color:rgb(228,247,251)}.S3aLQd .QkA63b:not(.RDPZE):hover,.S3aLQd .Y5sE8d:not(.RDPZE):hover,.S3aLQd .QkA63b:not(.RDPZE).u3bW4e,.S3aLQd .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(0,123,131,.2),0 1px 1px 0 rgba(0,123,131,.14),0 1px 3px 0 rgba(0,123,131,.12)}.S3aLQd .QkA63b:not(.RDPZE).iWO5td,.S3aLQd .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(0,123,131,.2),0 6px 10px 0 rgba(0,123,131,.14),0 1px 18px 0 rgba(0,123,131,.12)}.S3aLQd .DqwBN:not(.RDPZE),.S3aLQd .YhQJj:not(.RDPZE),.S3aLQd .K2V86d:not(.RDPZE),.S3aLQd .l3F1ye:not(.RDPZE),.S3aLQd .An19kf:not(.RDPZE),.S3aLQd .BEAGS:not(.RDPZE),.S3aLQd .AeAAkf:not(.RDPZE){color:rgb(0,123,131)}.S3aLQd .l3F1ye.j6PN2:not(.RDPZE){color:rgb(120,217,236)}.S3aLQd .wwnMtb:not(.RDPZE),.S3aLQd .OZ6W0d:not(.RDPZE){color:rgb(0,123,131);fill:rgb(0,123,131)}.S3aLQd .wwnMtb:not(.RDPZE):hover,.S3aLQd .OZ6W0d:not(.RDPZE):hover{background-color:rgba(0,123,131,.08)}.S3aLQd .wwnMtb:not(.RDPZE).u3bW4e,.S3aLQd .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(0,123,131,.12)}.S3aLQd .wwnMtb:not(.RDPZE).u3bW4e:hover,.S3aLQd .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(0,123,131,.16)}.S3aLQd .BEAGS.iWO5td,.S3aLQd .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(0,123,131,.2),0 1px 1px 0 rgba(0,123,131,.14),0 1px 3px 0 rgba(0,123,131,.12)}.S3aLQd .DqwBN .MbhUzd,.S3aLQd .YhQJj .MbhUzd,.S3aLQd .K2V86d .MbhUzd,.S3aLQd .l3F1ye .MbhUzd,.S3aLQd .BEAGS .MbhUzd,.S3aLQd .AeAAkf .MbhUzd,.S3aLQd .An19kf .MbhUzd,.S3aLQd .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(0,123,131,.16),rgba(0,123,131,.16) 80%,rgba(0,123,131,0) 100%)}.S3aLQd .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(120,217,236,.16),rgba(120,217,236,.16) 80%,rgba(120,217,236,0) 100%)}.S3aLQd .AeAAkf:not(.RDPZE) .CeoRYc,.S3aLQd .BEAGS:not(.RDPZE) .CeoRYc,.S3aLQd .An19kf:not(.RDPZE) .CeoRYc,.S3aLQd .l3F1ye:not(.RDPZE) .CeoRYc,.S3aLQd .YhQJj:not(.RDPZE) .CeoRYc,.S3aLQd .K2V86d:not(.RDPZE) .CeoRYc,.S3aLQd .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(0,123,131)}.S3aLQd .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(120,217,236)}.S3aLQd .AeAAkf:not(.RDPZE):hover,.S3aLQd .AeAAkf:not(.RDPZE).u3bW4e,.S3aLQd .BEAGS:not(.RDPZE):hover,.S3aLQd .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(18,158,175,.2)}.S3aLQd .DqwBN:not(.RDPZE):hover .CeoRYc,.S3aLQd .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.S3aLQd .YhQJj:not(.RDPZE):hover .CeoRYc,.S3aLQd .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.S3aLQd .K2V86d:not(.RDPZE):hover .CeoRYc,.S3aLQd .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.S3aLQd .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.S3aLQd .l3F1ye:not(.RDPZE):hover .CeoRYc,.S3aLQd .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(18,158,175)}.S3aLQd .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.S3aLQd .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(120,217,236)}.S3aLQd .aiSeRd:not(.RDPZE).N2RpBe,.S3aLQd .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(18,158,175)}.S3aLQd .aiSeRd:not(.RDPZE):hover .MbhUzd,.S3aLQd .aiSeRd:not(.RDPZE):focus .MbhUzd,.S3aLQd .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.S3aLQd .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(0,123,131,.08)}.S3aLQd .d7L4fc:hover .hYsg7c,.S3aLQd .NtlN8c:hover .hYsg7c{border-color:rgb(228,247,251)}.S3aLQd .d7L4fc:hover .MbhUzd,.S3aLQd .NtlN8c:hover .MbhUzd{background-color:rgba(0,123,131,.04)}.S3aLQd .d7L4fc .hYsg7c .nQOrEb,.S3aLQd .d7L4fc .hYsg7c.RDPZE .nQOrEb,.S3aLQd .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(18,158,175)}.S3aLQd .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.S3aLQd .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(0,123,131,.08)}.S3aLQd .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(18,158,175)}.S3aLQd .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#5ddfee}.S3aLQd .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(18,158,175,.3)}.S3aLQd .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#baf1f8}.S3aLQd .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(18,158,175,.04)}.S3aLQd .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.S3aLQd .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.S3aLQd .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(18,158,175,.12)}.S3aLQd .HyS0Qd:not(.RDPZE) .zHQkBf,.S3aLQd .fWf7qe:not(.RDPZE) .tL9Q4c,.S3aLQd .D3oBEe:not(.RDPZE) .zHQkBf,.S3aLQd .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(18,158,175)}.S3aLQd .HyS0Qd:not(.RDPZE) .cXrdqd,.S3aLQd .fWf7qe:not(.RDPZE) .cXrdqd,.S3aLQd .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(18,158,175)}.S3aLQd .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.S3aLQd .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(18,158,175)}.S3aLQd .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.S3aLQd .HyS0Qd input:not([disabled]):focus~.snByac,.S3aLQd .fWf7qe:not(.RDPZE).u3bW4e .snByac,.S3aLQd .D3oBEe:not(.RDPZE).u3bW4e .snByac,.S3aLQd .D3oBEe input:not([disabled]):focus~.snByac,.S3aLQd .AkVYk:not(.RDPZE).u3bW4e .snByac,.S3aLQd .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(0,123,131)}.S3aLQd .ybOdnf:not(.RDPZE).iWO5td,.S3aLQd .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.S3aLQd .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(228,247,251)}.S3aLQd .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(18,158,175);fill:rgb(18,158,175)}.S3aLQd .mRipsb{background-color:rgb(18,158,175)}.S3aLQd .bJuVn.KKjvXb{background-color:rgb(0,123,131)}.S3aLQd .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(0,123,131),transparent)}.S3aLQd .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(0,123,131),transparent)}.S3aLQd .bJuVn.u3bW4e.KKjvXb.KKjvXb,.S3aLQd .bJuVn.KKjvXb.KKjvXb:hover{background-color:#008d96}.S3aLQd .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.S3aLQd .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#008d96,transparent)}.S3aLQd .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.S3aLQd .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#008d96,transparent)}.S3aLQd .pAlOFe{color:rgb(0,123,131);fill:rgb(0,123,131)}.S3aLQd .bDxw8b:not(:disabled){background-color:rgb(0,123,131)}.S3aLQd .FL3Khc:not(:disabled){color:rgb(0,123,131)}.S3aLQd .FL3Khc:not(:disabled):hover{color:rgb(0,123,131)}.S3aLQd .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.S3aLQd .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(0,123,131)}.S3aLQd .FL3Khc .VfPpkd-Jh9lGc::before,.S3aLQd .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(0,123,131)}.S3aLQd .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.S3aLQd .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(0,123,131)}.S3aLQd .n42Gr:not(:disabled){color:rgb(0,123,131)}.S3aLQd .n42Gr:not(:disabled):hover{color:rgb(0,123,131)}.S3aLQd .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.S3aLQd .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(0,123,131)}.S3aLQd .n42Gr .VfPpkd-Jh9lGc::before,.S3aLQd .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(0,123,131)}.S3aLQd .J5y29e:not(:disabled){color:rgb(0,123,131)}.S3aLQd .J5y29e:not(:disabled):hover{color:rgb(0,123,131)}.S3aLQd .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.S3aLQd .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(0,123,131)}.S3aLQd .J5y29e .VfPpkd-Jh9lGc::before,.S3aLQd .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(0,123,131)}.S3aLQd .LgeCif{color:rgb(0,123,131)}.S3aLQd .LgeCif:disabled{color:rgba(60,64,67,.38)}.S3aLQd .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.S3aLQd .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(0,123,131)}.S3aLQd .wlZwYd:not(:disabled){background-color:rgb(228,247,251)}.S3aLQd .wlZwYd:not(:disabled){color:rgb(0,123,131)}.S3aLQd .wlZwYd:not(:disabled):hover{color:rgb(0,123,131)}.S3aLQd .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.S3aLQd .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(0,123,131)}.S3aLQd .wlZwYd .VfPpkd-Jh9lGc::before,.S3aLQd .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(0,123,131)}.S3aLQd .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.S3aLQd .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(18,158,175);border-color:var(--mdc-checkbox-selected-icon-color,rgb(18,158,175));background-color:rgb(18,158,175);background-color:var(--mdc-checkbox-selected-icon-color,rgb(18,158,175))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FF129EAF00000000FF129EAF{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(18,158,175);border-color:var(--mdc-checkbox-selected-icon-color,rgb(18,158,175));background-color:rgb(18,158,175);background-color:var(--mdc-checkbox-selected-icon-color,rgb(18,158,175))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FF129EAF00000000FF129EAF{0%,80%{border-color:rgb(18,158,175);border-color:var(--mdc-checkbox-selected-icon-color,rgb(18,158,175));background-color:rgb(18,158,175);background-color:var(--mdc-checkbox-selected-icon-color,rgb(18,158,175))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.S3aLQd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FF129EAF00000000FF129EAF}.S3aLQd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FF129EAF00000000FF129EAF}.S3aLQd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.S3aLQd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(0,123,131);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(0,123,131));background-color:rgb(0,123,131);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(0,123,131))}.S3aLQd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF007B8300000000FF007B83}.S3aLQd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF007B8300000000FF007B83}.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(0,123,131);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(0,123,131));background-color:rgb(0,123,131);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(0,123,131))}.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF007B8300000000FF007B83}.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF007B8300000000FF007B83}.S3aLQd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.S3aLQd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(0,123,131);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(0,123,131));background-color:rgb(0,123,131);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(0,123,131))}@keyframes mdc-checkbox-fade-in-background-FF202124FF007B8300000000FF007B83{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(0,123,131);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(0,123,131));background-color:rgb(0,123,131);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(0,123,131))}}@keyframes mdc-checkbox-fade-out-background-FF202124FF007B8300000000FF007B83{0%,80%{border-color:rgb(0,123,131);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(0,123,131));background-color:rgb(0,123,131);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(0,123,131))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.S3aLQd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF007B8300000000FF007B83}.S3aLQd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.S3aLQd .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF007B8300000000FF007B83}.S3aLQd .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.S3aLQd .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(0,123,131);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(0,123,131))}.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.S3aLQd .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(0,123,131);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(0,123,131))}.S3aLQd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.S3aLQd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.S3aLQd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.S3aLQd .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.S3aLQd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.S3aLQd .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(0,123,131)}.S3aLQd .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob:hover .VfPpkd-eHTEvd::before,.S3aLQd .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(0,123,131)}.S3aLQd .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(18,158,175)}.S3aLQd .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.S3aLQd .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(0,123,131)}.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(18,158,175)}.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(0,123,131)}.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(0,123,131)}.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(0,123,131)}.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(0,123,131)}.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(0,123,131)}.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.S3aLQd .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(0,123,131)}.S3aLQd .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#a1e3f1}.S3aLQd .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#a1e3f1}.S3aLQd .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#a1e3f1}.S3aLQd .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#a1e3f1}.S3aLQd .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(228,247,251)}.S3aLQd .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(0,123,131)}.S3aLQd .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(0,123,131)}.S3aLQd .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(0,123,131)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(18,158,175)}.S3aLQd .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.S3aLQd .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(18,158,175)}.S3aLQd .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.S3aLQd .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(18,158,175);background-color:var(--mdc-ripple-color,rgb(18,158,175))}.S3aLQd .U5B3me:not(:disabled){color:rgb(120,217,236)}.S3aLQd .U5B3me:not(:disabled):hover{color:rgb(120,217,236)}.S3aLQd .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.S3aLQd .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(120,217,236)}.S3aLQd .U5B3me .VfPpkd-Jh9lGc::before,.S3aLQd .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(120,217,236)}.S3aLQd .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(0,123,131)}.zvzLKc.bFjUmb-Ysl7Fe,.zvzLKc .bFjUmb-Ysl7Fe,.zvzLKc.CNpREd.bFjUmb-Ysl7Fe,.zvzLKc.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(253,231,243)}.zvzLKc.bFjUmb-Wvd9Cc,.zvzLKc .bFjUmb-Wvd9Cc,.zvzLKc.CNpREd.bFjUmb-Wvd9Cc,.zvzLKc.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(229,37,146)}.zvzLKc.bFjUmb-Tvm9db,.zvzLKc .bFjUmb-Tvm9db,.zvzLKc.CNpREd.bFjUmb-Tvm9db,.zvzLKc.CNpREd .bFjUmb-Tvm9db{background-color:rgb(184,6,114)}.zvzLKc.yxp05b-Wvd9Cc,.zvzLKc .yxp05b-Wvd9Cc,.zvzLKc.CNpREd.yxp05b-Wvd9Cc,.zvzLKc.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(229,37,146)}.zvzLKc.VnOHwf-Ysl7Fe,.zvzLKc .VnOHwf-Ysl7Fe,.zvzLKc.CNpREd.VnOHwf-Ysl7Fe,.zvzLKc.CNpREd .VnOHwf-Ysl7Fe{color:rgb(253,231,243);fill:rgb(253,231,243)}.zvzLKc.VnOHwf-Wvd9Cc,.zvzLKc .VnOHwf-Wvd9Cc,.zvzLKc.CNpREd.VnOHwf-Wvd9Cc,.zvzLKc.CNpREd .VnOHwf-Wvd9Cc{color:rgb(229,37,146);fill:rgb(229,37,146)}.zvzLKc.VnOHwf-Tvm9db,.zvzLKc .VnOHwf-Tvm9db,.zvzLKc.CNpREd.VnOHwf-Tvm9db,.zvzLKc.CNpREd .VnOHwf-Tvm9db{color:rgb(184,6,114);fill:rgb(184,6,114)}.zvzLKc.eL9Cfb,.zvzLKc .eL9Cfb,.zvzLKc.L5mE7d,.zvzLKc .L5mE7d,.zvzLKc.eL9Cfb:hover,.zvzLKc .eL9Cfb:hover,.zvzLKc.eL9Cfb:focus,.zvzLKc .eL9Cfb:focus,.zvzLKc.CNpREd.eL9Cfb,.zvzLKc.CNpREd .eL9Cfb,.zvzLKc.CNpREd.L5mE7d,.zvzLKc.CNpREd .L5mE7d,.zvzLKc.CNpREd.eL9Cfb:hover,.zvzLKc.CNpREd .eL9Cfb:hover,.zvzLKc.CNpREd.eL9Cfb:focus,.zvzLKc.CNpREd .eL9Cfb:focus{color:rgb(184,6,114)}.zvzLKc.L5mE7d:hover,.zvzLKc .L5mE7d:hover,.zvzLKc.L5mE7d:focus,.zvzLKc .L5mE7d:focus,.zvzLKc.L5mE7d:visited,.zvzLKc .L5mE7d:visited,.zvzLKc.CNpREd.L5mE7d:hover,.zvzLKc.CNpREd .L5mE7d:hover,.zvzLKc.CNpREd.L5mE7d:focus,.zvzLKc.CNpREd .L5mE7d:focus,.zvzLKc.CNpREd.L5mE7d:visited,.zvzLKc.CNpREd .L5mE7d:visited{color:rgb(229,37,146)}.zvzLKc .VUoKZ{background-color:rgb(253,231,243)}.zvzLKc .TRHLAc{background-color:rgb(229,37,146)}.zvzLKc .tgNIJf-Ysl7Fe:focus{border-color:rgb(253,231,243)}.zvzLKc .cjzpkc-Wvd9Cc:focus-within,.zvzLKc .tgNIJf-Wvd9Cc:focus{border-color:rgb(229,37,146)}.zvzLKc .u3bW4e .zZN2Lb-Wvd9Cc,.zvzLKc .zZN2Lb-Wvd9Cc:focus,.zvzLKc .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(229,37,146)}.zvzLKc .P3W0Dd-Ysl7Fe:focus,.zvzLKc.maXJsd:focus .P3W0Dd-Ysl7Fe,.zvzLKc .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(253,231,243)}.zvzLKc .VBEdtc-Wvd9Cc:hover,.zvzLKc.MymH0d:hover .VBEdtc-Wvd9Cc,.zvzLKc .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(229,37,146)}.zvzLKc.MymH0d:hover .UISY8d-Tvm9db,.zvzLKc.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.zvzLKc .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(229,37,146)}.zvzLKc .UISY8d-Ysl7Fe:hover,.zvzLKc.MymH0d:hover .UISY8d-Ysl7Fe,.zvzLKc .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(253,231,243)}.zvzLKc .mxmXhf{color:rgb(184,6,114);fill:rgb(184,6,114)}.zvzLKc .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.zvzLKc .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.zvzLKc .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.zvzLKc .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.zvzLKc .ZoT1D:focus-within.boxOzd,.zvzLKc .ZoT1D:focus-within.idtp4e,.zvzLKc .ZoT1D :focus-within.boxOzd,.zvzLKc .ZoT1D :focus-within.idtp4e{background-color:rgb(253,231,243)}.zvzLKc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.zvzLKc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.zvzLKc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.zvzLKc .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.zvzLKc .ZoT1D:hover.j6KDAd,.zvzLKc .ZoT1D:hover.idtp4e,.zvzLKc .ZoT1D:hover .j6KDAd,.zvzLKc .ZoT1D:hover .idtp4e{background-color:rgb(253,231,243)}.zvzLKc .OGhwGf:hover,.zvzLKc .OGhwGf:focus{color:rgb(184,6,114)}.zvzLKc .ra2NV,.zvzLKc.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(229,37,146),transparent)}.zvzLKc .eumXzf:after{border-color:rgb(184,6,114)}.zvzLKc .zKHdkd .cXrdqd,.zvzLKc .kPBwDb{background-color:rgb(229,37,146)}.zvzLKc .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.zvzLKc .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(229,37,146)}.zvzLKc .bkIpNd .uHMk6b{border-color:rgb(253,231,243)}.zvzLKc .zJKIV .nQOrEb,.zvzLKc .zJKIV.RDPZE .nQOrEb,.zvzLKc .zJKIV.N2RpBe .Id5V1,.zvzLKc .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(229,37,146)}.zvzLKc .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(229,37,146);opacity:.5}.zvzLKc .zJKIV.i9xfbb>.MbhUzd,.zvzLKc .zJKIV.u3bW4e>.MbhUzd,.zvzLKc .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.zvzLKc .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(253,231,243)}.zvzLKc .HQ8yf:not(.RDPZE),.zvzLKc .HQ8yf:not(.RDPZE) a{color:rgb(229,37,146)}.zvzLKc .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(229,37,146,.15)}.zvzLKc .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(229,37,146,.25),rgba(229,37,146,.25) 80%,rgb(229,37,146) 100%)}.zvzLKc .uO32ac,.zvzLKc .ypv4re{border-bottom:1px solid rgb(229,37,146)}.zvzLKc .DqwBN:not(.RDPZE) .TpQm9d,.zvzLKc .l3F1ye:not(.RDPZE) .TpQm9d,.zvzLKc .YhQJj:not(.RDPZE) .TpQm9d,.zvzLKc .K2V86d:not(.RDPZE) .TpQm9d,.zvzLKc .An19kf:not(.RDPZE) .TpQm9d{color:rgb(184,6,114);fill:rgb(184,6,114)}.zvzLKc .DqwBN .TpQm9d,.zvzLKc .YhQJj .TpQm9d,.zvzLKc .K2V86d .TpQm9d,.zvzLKc .l3F1ye .TpQm9d,.zvzLKc .An19kf .TpQm9d{color:rgb(184,6,114);fill:rgb(184,6,114)}.zvzLKc .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(255,139,203);fill:rgb(255,139,203)}.zvzLKc .QkA63b:not(.RDPZE),.zvzLKc .Y5sE8d:not(.RDPZE){background-color:rgb(184,6,114)}.zvzLKc .An19kf:not(.RDPZE){background-color:rgb(253,231,243)}.zvzLKc .QkA63b:not(.RDPZE):hover,.zvzLKc .Y5sE8d:not(.RDPZE):hover,.zvzLKc .QkA63b:not(.RDPZE).u3bW4e,.zvzLKc .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(184,6,114,.2),0 1px 1px 0 rgba(184,6,114,.14),0 1px 3px 0 rgba(184,6,114,.12)}.zvzLKc .QkA63b:not(.RDPZE).iWO5td,.zvzLKc .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(184,6,114,.2),0 6px 10px 0 rgba(184,6,114,.14),0 1px 18px 0 rgba(184,6,114,.12)}.zvzLKc .DqwBN:not(.RDPZE),.zvzLKc .YhQJj:not(.RDPZE),.zvzLKc .K2V86d:not(.RDPZE),.zvzLKc .l3F1ye:not(.RDPZE),.zvzLKc .An19kf:not(.RDPZE),.zvzLKc .BEAGS:not(.RDPZE),.zvzLKc .AeAAkf:not(.RDPZE){color:rgb(184,6,114)}.zvzLKc .l3F1ye.j6PN2:not(.RDPZE){color:rgb(255,139,203)}.zvzLKc .wwnMtb:not(.RDPZE),.zvzLKc .OZ6W0d:not(.RDPZE){color:rgb(184,6,114);fill:rgb(184,6,114)}.zvzLKc .wwnMtb:not(.RDPZE):hover,.zvzLKc .OZ6W0d:not(.RDPZE):hover{background-color:rgba(184,6,114,.08)}.zvzLKc .wwnMtb:not(.RDPZE).u3bW4e,.zvzLKc .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(184,6,114,.12)}.zvzLKc .wwnMtb:not(.RDPZE).u3bW4e:hover,.zvzLKc .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(184,6,114,.16)}.zvzLKc .BEAGS.iWO5td,.zvzLKc .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(184,6,114,.2),0 1px 1px 0 rgba(184,6,114,.14),0 1px 3px 0 rgba(184,6,114,.12)}.zvzLKc .DqwBN .MbhUzd,.zvzLKc .YhQJj .MbhUzd,.zvzLKc .K2V86d .MbhUzd,.zvzLKc .l3F1ye .MbhUzd,.zvzLKc .BEAGS .MbhUzd,.zvzLKc .AeAAkf .MbhUzd,.zvzLKc .An19kf .MbhUzd,.zvzLKc .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(184,6,114,.16),rgba(184,6,114,.16) 80%,rgba(184,6,114,0) 100%)}.zvzLKc .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(255,139,203,.16),rgba(255,139,203,.16) 80%,rgba(255,139,203,0) 100%)}.zvzLKc .AeAAkf:not(.RDPZE) .CeoRYc,.zvzLKc .BEAGS:not(.RDPZE) .CeoRYc,.zvzLKc .An19kf:not(.RDPZE) .CeoRYc,.zvzLKc .l3F1ye:not(.RDPZE) .CeoRYc,.zvzLKc .YhQJj:not(.RDPZE) .CeoRYc,.zvzLKc .K2V86d:not(.RDPZE) .CeoRYc,.zvzLKc .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(184,6,114)}.zvzLKc .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(255,139,203)}.zvzLKc .AeAAkf:not(.RDPZE):hover,.zvzLKc .AeAAkf:not(.RDPZE).u3bW4e,.zvzLKc .BEAGS:not(.RDPZE):hover,.zvzLKc .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(229,37,146,.2)}.zvzLKc .DqwBN:not(.RDPZE):hover .CeoRYc,.zvzLKc .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.zvzLKc .YhQJj:not(.RDPZE):hover .CeoRYc,.zvzLKc .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.zvzLKc .K2V86d:not(.RDPZE):hover .CeoRYc,.zvzLKc .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.zvzLKc .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.zvzLKc .l3F1ye:not(.RDPZE):hover .CeoRYc,.zvzLKc .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(229,37,146)}.zvzLKc .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.zvzLKc .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(255,139,203)}.zvzLKc .aiSeRd:not(.RDPZE).N2RpBe,.zvzLKc .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(229,37,146)}.zvzLKc .aiSeRd:not(.RDPZE):hover .MbhUzd,.zvzLKc .aiSeRd:not(.RDPZE):focus .MbhUzd,.zvzLKc .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.zvzLKc .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(184,6,114,.08)}.zvzLKc .d7L4fc:hover .hYsg7c,.zvzLKc .NtlN8c:hover .hYsg7c{border-color:rgb(253,231,243)}.zvzLKc .d7L4fc:hover .MbhUzd,.zvzLKc .NtlN8c:hover .MbhUzd{background-color:rgba(184,6,114,.04)}.zvzLKc .d7L4fc .hYsg7c .nQOrEb,.zvzLKc .d7L4fc .hYsg7c.RDPZE .nQOrEb,.zvzLKc .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(229,37,146)}.zvzLKc .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.zvzLKc .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(184,6,114,.08)}.zvzLKc .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(229,37,146)}.zvzLKc .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#ec60af}.zvzLKc .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(229,37,146,.3)}.zvzLKc .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#f7bbdd}.zvzLKc .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(229,37,146,.04)}.zvzLKc .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.zvzLKc .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.zvzLKc .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(229,37,146,.12)}.zvzLKc .HyS0Qd:not(.RDPZE) .zHQkBf,.zvzLKc .fWf7qe:not(.RDPZE) .tL9Q4c,.zvzLKc .D3oBEe:not(.RDPZE) .zHQkBf,.zvzLKc .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(229,37,146)}.zvzLKc .HyS0Qd:not(.RDPZE) .cXrdqd,.zvzLKc .fWf7qe:not(.RDPZE) .cXrdqd,.zvzLKc .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(229,37,146)}.zvzLKc .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.zvzLKc .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(229,37,146)}.zvzLKc .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.zvzLKc .HyS0Qd input:not([disabled]):focus~.snByac,.zvzLKc .fWf7qe:not(.RDPZE).u3bW4e .snByac,.zvzLKc .D3oBEe:not(.RDPZE).u3bW4e .snByac,.zvzLKc .D3oBEe input:not([disabled]):focus~.snByac,.zvzLKc .AkVYk:not(.RDPZE).u3bW4e .snByac,.zvzLKc .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(184,6,114)}.zvzLKc .ybOdnf:not(.RDPZE).iWO5td,.zvzLKc .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.zvzLKc .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(253,231,243)}.zvzLKc .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(229,37,146);fill:rgb(229,37,146)}.zvzLKc .mRipsb{background-color:rgb(229,37,146)}.zvzLKc .bJuVn.KKjvXb{background-color:rgb(184,6,114)}.zvzLKc .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(184,6,114),transparent)}.zvzLKc .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(184,6,114),transparent)}.zvzLKc .bJuVn.u3bW4e.KKjvXb.KKjvXb,.zvzLKc .bJuVn.KKjvXb.KKjvXb:hover{background-color:#c7077c}.zvzLKc .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.zvzLKc .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#c7077c,transparent)}.zvzLKc .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.zvzLKc .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#c7077c,transparent)}.zvzLKc .pAlOFe{color:rgb(184,6,114);fill:rgb(184,6,114)}.zvzLKc .bDxw8b:not(:disabled){background-color:rgb(184,6,114)}.zvzLKc .FL3Khc:not(:disabled){color:rgb(184,6,114)}.zvzLKc .FL3Khc:not(:disabled):hover{color:rgb(184,6,114)}.zvzLKc .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.zvzLKc .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(184,6,114)}.zvzLKc .FL3Khc .VfPpkd-Jh9lGc::before,.zvzLKc .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(184,6,114)}.zvzLKc .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.zvzLKc .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(184,6,114)}.zvzLKc .n42Gr:not(:disabled){color:rgb(184,6,114)}.zvzLKc .n42Gr:not(:disabled):hover{color:rgb(184,6,114)}.zvzLKc .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.zvzLKc .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(184,6,114)}.zvzLKc .n42Gr .VfPpkd-Jh9lGc::before,.zvzLKc .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(184,6,114)}.zvzLKc .J5y29e:not(:disabled){color:rgb(184,6,114)}.zvzLKc .J5y29e:not(:disabled):hover{color:rgb(184,6,114)}.zvzLKc .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.zvzLKc .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(184,6,114)}.zvzLKc .J5y29e .VfPpkd-Jh9lGc::before,.zvzLKc .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(184,6,114)}.zvzLKc .LgeCif{color:rgb(184,6,114)}.zvzLKc .LgeCif:disabled{color:rgba(60,64,67,.38)}.zvzLKc .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.zvzLKc .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(184,6,114)}.zvzLKc .wlZwYd:not(:disabled){background-color:rgb(253,231,243)}.zvzLKc .wlZwYd:not(:disabled){color:rgb(184,6,114)}.zvzLKc .wlZwYd:not(:disabled):hover{color:rgb(184,6,114)}.zvzLKc .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.zvzLKc .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(184,6,114)}.zvzLKc .wlZwYd .VfPpkd-Jh9lGc::before,.zvzLKc .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(184,6,114)}.zvzLKc .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.zvzLKc .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(229,37,146);border-color:var(--mdc-checkbox-selected-icon-color,rgb(229,37,146));background-color:rgb(229,37,146);background-color:var(--mdc-checkbox-selected-icon-color,rgb(229,37,146))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FFE5259200000000FFE52592{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(229,37,146);border-color:var(--mdc-checkbox-selected-icon-color,rgb(229,37,146));background-color:rgb(229,37,146);background-color:var(--mdc-checkbox-selected-icon-color,rgb(229,37,146))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FFE5259200000000FFE52592{0%,80%{border-color:rgb(229,37,146);border-color:var(--mdc-checkbox-selected-icon-color,rgb(229,37,146));background-color:rgb(229,37,146);background-color:var(--mdc-checkbox-selected-icon-color,rgb(229,37,146))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.zvzLKc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FFE5259200000000FFE52592}.zvzLKc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FFE5259200000000FFE52592}.zvzLKc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.zvzLKc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(184,6,114);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(184,6,114));background-color:rgb(184,6,114);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(184,6,114))}.zvzLKc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FFB8067200000000FFB80672}.zvzLKc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FFB8067200000000FFB80672}.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(184,6,114);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(184,6,114));background-color:rgb(184,6,114);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(184,6,114))}.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FFB8067200000000FFB80672}.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FFB8067200000000FFB80672}.zvzLKc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.zvzLKc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(184,6,114);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(184,6,114));background-color:rgb(184,6,114);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(184,6,114))}@keyframes mdc-checkbox-fade-in-background-FF202124FFB8067200000000FFB80672{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(184,6,114);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(184,6,114));background-color:rgb(184,6,114);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(184,6,114))}}@keyframes mdc-checkbox-fade-out-background-FF202124FFB8067200000000FFB80672{0%,80%{border-color:rgb(184,6,114);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(184,6,114));background-color:rgb(184,6,114);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(184,6,114))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.zvzLKc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FFB8067200000000FFB80672}.zvzLKc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.zvzLKc .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FFB8067200000000FFB80672}.zvzLKc .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.zvzLKc .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(184,6,114);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(184,6,114))}.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.zvzLKc .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(184,6,114);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(184,6,114))}.zvzLKc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.zvzLKc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.zvzLKc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.zvzLKc .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.zvzLKc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.zvzLKc .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(184,6,114)}.zvzLKc .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob:hover .VfPpkd-eHTEvd::before,.zvzLKc .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(184,6,114)}.zvzLKc .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(229,37,146)}.zvzLKc .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.zvzLKc .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(184,6,114)}.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(229,37,146)}.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(184,6,114)}.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(184,6,114)}.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(184,6,114)}.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(184,6,114)}.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(184,6,114)}.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.zvzLKc .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(184,6,114)}.zvzLKc .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#f7a0d0}.zvzLKc .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#f7a0d0}.zvzLKc .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#f7a0d0}.zvzLKc .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#f7a0d0}.zvzLKc .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(253,231,243)}.zvzLKc .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(184,6,114)}.zvzLKc .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(184,6,114)}.zvzLKc .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(184,6,114)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(229,37,146)}.zvzLKc .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.zvzLKc .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(229,37,146)}.zvzLKc .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.zvzLKc .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(229,37,146);background-color:var(--mdc-ripple-color,rgb(229,37,146))}.zvzLKc .U5B3me:not(:disabled){color:rgb(255,139,203)}.zvzLKc .U5B3me:not(:disabled):hover{color:rgb(255,139,203)}.zvzLKc .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.zvzLKc .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(255,139,203)}.zvzLKc .U5B3me .VfPpkd-Jh9lGc::before,.zvzLKc .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(255,139,203)}.zvzLKc .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(184,6,114)}.WFUiUb.bFjUmb-Ysl7Fe,.WFUiUb .bFjUmb-Ysl7Fe,.WFUiUb.CNpREd.bFjUmb-Ysl7Fe,.WFUiUb.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(230,244,234)}.WFUiUb.bFjUmb-Wvd9Cc,.WFUiUb .bFjUmb-Wvd9Cc,.WFUiUb.CNpREd.bFjUmb-Wvd9Cc,.WFUiUb.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(30,142,62)}.WFUiUb.bFjUmb-Tvm9db,.WFUiUb .bFjUmb-Tvm9db,.WFUiUb.CNpREd.bFjUmb-Tvm9db,.WFUiUb.CNpREd .bFjUmb-Tvm9db{background-color:rgb(19,115,51)}.WFUiUb.yxp05b-Wvd9Cc,.WFUiUb .yxp05b-Wvd9Cc,.WFUiUb.CNpREd.yxp05b-Wvd9Cc,.WFUiUb.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(30,142,62)}.WFUiUb.VnOHwf-Ysl7Fe,.WFUiUb .VnOHwf-Ysl7Fe,.WFUiUb.CNpREd.VnOHwf-Ysl7Fe,.WFUiUb.CNpREd .VnOHwf-Ysl7Fe{color:rgb(230,244,234);fill:rgb(230,244,234)}.WFUiUb.VnOHwf-Wvd9Cc,.WFUiUb .VnOHwf-Wvd9Cc,.WFUiUb.CNpREd.VnOHwf-Wvd9Cc,.WFUiUb.CNpREd .VnOHwf-Wvd9Cc{color:rgb(30,142,62);fill:rgb(30,142,62)}.WFUiUb.VnOHwf-Tvm9db,.WFUiUb .VnOHwf-Tvm9db,.WFUiUb.CNpREd.VnOHwf-Tvm9db,.WFUiUb.CNpREd .VnOHwf-Tvm9db{color:rgb(19,115,51);fill:rgb(19,115,51)}.WFUiUb.eL9Cfb,.WFUiUb .eL9Cfb,.WFUiUb.L5mE7d,.WFUiUb .L5mE7d,.WFUiUb.eL9Cfb:hover,.WFUiUb .eL9Cfb:hover,.WFUiUb.eL9Cfb:focus,.WFUiUb .eL9Cfb:focus,.WFUiUb.CNpREd.eL9Cfb,.WFUiUb.CNpREd .eL9Cfb,.WFUiUb.CNpREd.L5mE7d,.WFUiUb.CNpREd .L5mE7d,.WFUiUb.CNpREd.eL9Cfb:hover,.WFUiUb.CNpREd .eL9Cfb:hover,.WFUiUb.CNpREd.eL9Cfb:focus,.WFUiUb.CNpREd .eL9Cfb:focus{color:rgb(19,115,51)}.WFUiUb.L5mE7d:hover,.WFUiUb .L5mE7d:hover,.WFUiUb.L5mE7d:focus,.WFUiUb .L5mE7d:focus,.WFUiUb.L5mE7d:visited,.WFUiUb .L5mE7d:visited,.WFUiUb.CNpREd.L5mE7d:hover,.WFUiUb.CNpREd .L5mE7d:hover,.WFUiUb.CNpREd.L5mE7d:focus,.WFUiUb.CNpREd .L5mE7d:focus,.WFUiUb.CNpREd.L5mE7d:visited,.WFUiUb.CNpREd .L5mE7d:visited{color:rgb(30,142,62)}.WFUiUb .VUoKZ{background-color:rgb(230,244,234)}.WFUiUb .TRHLAc{background-color:rgb(30,142,62)}.WFUiUb .tgNIJf-Ysl7Fe:focus{border-color:rgb(230,244,234)}.WFUiUb .cjzpkc-Wvd9Cc:focus-within,.WFUiUb .tgNIJf-Wvd9Cc:focus{border-color:rgb(30,142,62)}.WFUiUb .u3bW4e .zZN2Lb-Wvd9Cc,.WFUiUb .zZN2Lb-Wvd9Cc:focus,.WFUiUb .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(30,142,62)}.WFUiUb .P3W0Dd-Ysl7Fe:focus,.WFUiUb.maXJsd:focus .P3W0Dd-Ysl7Fe,.WFUiUb .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(230,244,234)}.WFUiUb .VBEdtc-Wvd9Cc:hover,.WFUiUb.MymH0d:hover .VBEdtc-Wvd9Cc,.WFUiUb .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(30,142,62)}.WFUiUb.MymH0d:hover .UISY8d-Tvm9db,.WFUiUb.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.WFUiUb .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(30,142,62)}.WFUiUb .UISY8d-Ysl7Fe:hover,.WFUiUb.MymH0d:hover .UISY8d-Ysl7Fe,.WFUiUb .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(230,244,234)}.WFUiUb .mxmXhf{color:rgb(19,115,51);fill:rgb(19,115,51)}.WFUiUb .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.WFUiUb .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.WFUiUb .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.WFUiUb .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.WFUiUb .ZoT1D:focus-within.boxOzd,.WFUiUb .ZoT1D:focus-within.idtp4e,.WFUiUb .ZoT1D :focus-within.boxOzd,.WFUiUb .ZoT1D :focus-within.idtp4e{background-color:rgb(230,244,234)}.WFUiUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.WFUiUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.WFUiUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.WFUiUb .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.WFUiUb .ZoT1D:hover.j6KDAd,.WFUiUb .ZoT1D:hover.idtp4e,.WFUiUb .ZoT1D:hover .j6KDAd,.WFUiUb .ZoT1D:hover .idtp4e{background-color:rgb(230,244,234)}.WFUiUb .OGhwGf:hover,.WFUiUb .OGhwGf:focus{color:rgb(19,115,51)}.WFUiUb .ra2NV,.WFUiUb.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(30,142,62),transparent)}.WFUiUb .eumXzf:after{border-color:rgb(19,115,51)}.WFUiUb .zKHdkd .cXrdqd,.WFUiUb .kPBwDb{background-color:rgb(30,142,62)}.WFUiUb .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.WFUiUb .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(30,142,62)}.WFUiUb .bkIpNd .uHMk6b{border-color:rgb(230,244,234)}.WFUiUb .zJKIV .nQOrEb,.WFUiUb .zJKIV.RDPZE .nQOrEb,.WFUiUb .zJKIV.N2RpBe .Id5V1,.WFUiUb .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(30,142,62)}.WFUiUb .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(30,142,62);opacity:.5}.WFUiUb .zJKIV.i9xfbb>.MbhUzd,.WFUiUb .zJKIV.u3bW4e>.MbhUzd,.WFUiUb .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.WFUiUb .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(230,244,234)}.WFUiUb .HQ8yf:not(.RDPZE),.WFUiUb .HQ8yf:not(.RDPZE) a{color:rgb(30,142,62)}.WFUiUb .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(30,142,62,.15)}.WFUiUb .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(30,142,62,.25),rgba(30,142,62,.25) 80%,rgb(30,142,62) 100%)}.WFUiUb .uO32ac,.WFUiUb .ypv4re{border-bottom:1px solid rgb(30,142,62)}.WFUiUb .DqwBN:not(.RDPZE) .TpQm9d,.WFUiUb .l3F1ye:not(.RDPZE) .TpQm9d,.WFUiUb .YhQJj:not(.RDPZE) .TpQm9d,.WFUiUb .K2V86d:not(.RDPZE) .TpQm9d,.WFUiUb .An19kf:not(.RDPZE) .TpQm9d{color:rgb(19,115,51);fill:rgb(19,115,51)}.WFUiUb .DqwBN .TpQm9d,.WFUiUb .YhQJj .TpQm9d,.WFUiUb .K2V86d .TpQm9d,.WFUiUb .l3F1ye .TpQm9d,.WFUiUb .An19kf .TpQm9d{color:rgb(19,115,51);fill:rgb(19,115,51)}.WFUiUb .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(129,201,149);fill:rgb(129,201,149)}.WFUiUb .QkA63b:not(.RDPZE),.WFUiUb .Y5sE8d:not(.RDPZE){background-color:rgb(19,115,51)}.WFUiUb .An19kf:not(.RDPZE){background-color:rgb(230,244,234)}.WFUiUb .QkA63b:not(.RDPZE):hover,.WFUiUb .Y5sE8d:not(.RDPZE):hover,.WFUiUb .QkA63b:not(.RDPZE).u3bW4e,.WFUiUb .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(19,115,51,.2),0 1px 1px 0 rgba(19,115,51,.14),0 1px 3px 0 rgba(19,115,51,.12)}.WFUiUb .QkA63b:not(.RDPZE).iWO5td,.WFUiUb .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(19,115,51,.2),0 6px 10px 0 rgba(19,115,51,.14),0 1px 18px 0 rgba(19,115,51,.12)}.WFUiUb .DqwBN:not(.RDPZE),.WFUiUb .YhQJj:not(.RDPZE),.WFUiUb .K2V86d:not(.RDPZE),.WFUiUb .l3F1ye:not(.RDPZE),.WFUiUb .An19kf:not(.RDPZE),.WFUiUb .BEAGS:not(.RDPZE),.WFUiUb .AeAAkf:not(.RDPZE){color:rgb(19,115,51)}.WFUiUb .l3F1ye.j6PN2:not(.RDPZE){color:rgb(129,201,149)}.WFUiUb .wwnMtb:not(.RDPZE),.WFUiUb .OZ6W0d:not(.RDPZE){color:rgb(19,115,51);fill:rgb(19,115,51)}.WFUiUb .wwnMtb:not(.RDPZE):hover,.WFUiUb .OZ6W0d:not(.RDPZE):hover{background-color:rgba(19,115,51,.08)}.WFUiUb .wwnMtb:not(.RDPZE).u3bW4e,.WFUiUb .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(19,115,51,.12)}.WFUiUb .wwnMtb:not(.RDPZE).u3bW4e:hover,.WFUiUb .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(19,115,51,.16)}.WFUiUb .BEAGS.iWO5td,.WFUiUb .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(19,115,51,.2),0 1px 1px 0 rgba(19,115,51,.14),0 1px 3px 0 rgba(19,115,51,.12)}.WFUiUb .DqwBN .MbhUzd,.WFUiUb .YhQJj .MbhUzd,.WFUiUb .K2V86d .MbhUzd,.WFUiUb .l3F1ye .MbhUzd,.WFUiUb .BEAGS .MbhUzd,.WFUiUb .AeAAkf .MbhUzd,.WFUiUb .An19kf .MbhUzd,.WFUiUb .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(19,115,51,.16),rgba(19,115,51,.16) 80%,rgba(19,115,51,0) 100%)}.WFUiUb .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(129,201,149,.16),rgba(129,201,149,.16) 80%,rgba(129,201,149,0) 100%)}.WFUiUb .AeAAkf:not(.RDPZE) .CeoRYc,.WFUiUb .BEAGS:not(.RDPZE) .CeoRYc,.WFUiUb .An19kf:not(.RDPZE) .CeoRYc,.WFUiUb .l3F1ye:not(.RDPZE) .CeoRYc,.WFUiUb .YhQJj:not(.RDPZE) .CeoRYc,.WFUiUb .K2V86d:not(.RDPZE) .CeoRYc,.WFUiUb .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(19,115,51)}.WFUiUb .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(129,201,149)}.WFUiUb .AeAAkf:not(.RDPZE):hover,.WFUiUb .AeAAkf:not(.RDPZE).u3bW4e,.WFUiUb .BEAGS:not(.RDPZE):hover,.WFUiUb .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(30,142,62,.2)}.WFUiUb .DqwBN:not(.RDPZE):hover .CeoRYc,.WFUiUb .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.WFUiUb .YhQJj:not(.RDPZE):hover .CeoRYc,.WFUiUb .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.WFUiUb .K2V86d:not(.RDPZE):hover .CeoRYc,.WFUiUb .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.WFUiUb .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.WFUiUb .l3F1ye:not(.RDPZE):hover .CeoRYc,.WFUiUb .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(30,142,62)}.WFUiUb .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.WFUiUb .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(129,201,149)}.WFUiUb .aiSeRd:not(.RDPZE).N2RpBe,.WFUiUb .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(30,142,62)}.WFUiUb .aiSeRd:not(.RDPZE):hover .MbhUzd,.WFUiUb .aiSeRd:not(.RDPZE):focus .MbhUzd,.WFUiUb .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.WFUiUb .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(19,115,51,.08)}.WFUiUb .d7L4fc:hover .hYsg7c,.WFUiUb .NtlN8c:hover .hYsg7c{border-color:rgb(230,244,234)}.WFUiUb .d7L4fc:hover .MbhUzd,.WFUiUb .NtlN8c:hover .MbhUzd{background-color:rgba(19,115,51,.04)}.WFUiUb .d7L4fc .hYsg7c .nQOrEb,.WFUiUb .d7L4fc .hYsg7c.RDPZE .nQOrEb,.WFUiUb .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(30,142,62)}.WFUiUb .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.WFUiUb .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(19,115,51,.08)}.WFUiUb .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(30,142,62)}.WFUiUb .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#6ce08d}.WFUiUb .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(30,142,62,.3)}.WFUiUb .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#c0f2ce}.WFUiUb .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(30,142,62,.04)}.WFUiUb .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.WFUiUb .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.WFUiUb .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(30,142,62,.12)}.WFUiUb .HyS0Qd:not(.RDPZE) .zHQkBf,.WFUiUb .fWf7qe:not(.RDPZE) .tL9Q4c,.WFUiUb .D3oBEe:not(.RDPZE) .zHQkBf,.WFUiUb .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(30,142,62)}.WFUiUb .HyS0Qd:not(.RDPZE) .cXrdqd,.WFUiUb .fWf7qe:not(.RDPZE) .cXrdqd,.WFUiUb .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(30,142,62)}.WFUiUb .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.WFUiUb .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(30,142,62)}.WFUiUb .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.WFUiUb .HyS0Qd input:not([disabled]):focus~.snByac,.WFUiUb .fWf7qe:not(.RDPZE).u3bW4e .snByac,.WFUiUb .D3oBEe:not(.RDPZE).u3bW4e .snByac,.WFUiUb .D3oBEe input:not([disabled]):focus~.snByac,.WFUiUb .AkVYk:not(.RDPZE).u3bW4e .snByac,.WFUiUb .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(19,115,51)}.WFUiUb .ybOdnf:not(.RDPZE).iWO5td,.WFUiUb .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.WFUiUb .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(230,244,234)}.WFUiUb .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(30,142,62);fill:rgb(30,142,62)}.WFUiUb .mRipsb{background-color:rgb(30,142,62)}.WFUiUb .bJuVn.KKjvXb{background-color:rgb(19,115,51)}.WFUiUb .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(19,115,51),transparent)}.WFUiUb .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(19,115,51),transparent)}.WFUiUb .bJuVn.u3bW4e.KKjvXb.KKjvXb,.WFUiUb .bJuVn.KKjvXb.KKjvXb:hover{background-color:#16833a}.WFUiUb .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.WFUiUb .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#16833a,transparent)}.WFUiUb .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.WFUiUb .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#16833a,transparent)}.WFUiUb .pAlOFe{color:rgb(19,115,51);fill:rgb(19,115,51)}.WFUiUb .bDxw8b:not(:disabled){background-color:rgb(19,115,51)}.WFUiUb .FL3Khc:not(:disabled){color:rgb(19,115,51)}.WFUiUb .FL3Khc:not(:disabled):hover{color:rgb(19,115,51)}.WFUiUb .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.WFUiUb .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(19,115,51)}.WFUiUb .FL3Khc .VfPpkd-Jh9lGc::before,.WFUiUb .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(19,115,51)}.WFUiUb .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.WFUiUb .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(19,115,51)}.WFUiUb .n42Gr:not(:disabled){color:rgb(19,115,51)}.WFUiUb .n42Gr:not(:disabled):hover{color:rgb(19,115,51)}.WFUiUb .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.WFUiUb .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(19,115,51)}.WFUiUb .n42Gr .VfPpkd-Jh9lGc::before,.WFUiUb .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(19,115,51)}.WFUiUb .J5y29e:not(:disabled){color:rgb(19,115,51)}.WFUiUb .J5y29e:not(:disabled):hover{color:rgb(19,115,51)}.WFUiUb .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.WFUiUb .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(19,115,51)}.WFUiUb .J5y29e .VfPpkd-Jh9lGc::before,.WFUiUb .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(19,115,51)}.WFUiUb .LgeCif{color:rgb(19,115,51)}.WFUiUb .LgeCif:disabled{color:rgba(60,64,67,.38)}.WFUiUb .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.WFUiUb .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(19,115,51)}.WFUiUb .wlZwYd:not(:disabled){background-color:rgb(230,244,234)}.WFUiUb .wlZwYd:not(:disabled){color:rgb(19,115,51)}.WFUiUb .wlZwYd:not(:disabled):hover{color:rgb(19,115,51)}.WFUiUb .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.WFUiUb .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(19,115,51)}.WFUiUb .wlZwYd .VfPpkd-Jh9lGc::before,.WFUiUb .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(19,115,51)}.WFUiUb .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.WFUiUb .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(30,142,62);border-color:var(--mdc-checkbox-selected-icon-color,rgb(30,142,62));background-color:rgb(30,142,62);background-color:var(--mdc-checkbox-selected-icon-color,rgb(30,142,62))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FF1E8E3E00000000FF1E8E3E{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(30,142,62);border-color:var(--mdc-checkbox-selected-icon-color,rgb(30,142,62));background-color:rgb(30,142,62);background-color:var(--mdc-checkbox-selected-icon-color,rgb(30,142,62))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FF1E8E3E00000000FF1E8E3E{0%,80%{border-color:rgb(30,142,62);border-color:var(--mdc-checkbox-selected-icon-color,rgb(30,142,62));background-color:rgb(30,142,62);background-color:var(--mdc-checkbox-selected-icon-color,rgb(30,142,62))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.WFUiUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FF1E8E3E00000000FF1E8E3E}.WFUiUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FF1E8E3E00000000FF1E8E3E}.WFUiUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.WFUiUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(19,115,51);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(19,115,51));background-color:rgb(19,115,51);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(19,115,51))}.WFUiUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF13733300000000FF137333}.WFUiUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF13733300000000FF137333}.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(19,115,51);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(19,115,51));background-color:rgb(19,115,51);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(19,115,51))}.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF13733300000000FF137333}.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF13733300000000FF137333}.WFUiUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.WFUiUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(19,115,51);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(19,115,51));background-color:rgb(19,115,51);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(19,115,51))}@keyframes mdc-checkbox-fade-in-background-FF202124FF13733300000000FF137333{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(19,115,51);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(19,115,51));background-color:rgb(19,115,51);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(19,115,51))}}@keyframes mdc-checkbox-fade-out-background-FF202124FF13733300000000FF137333{0%,80%{border-color:rgb(19,115,51);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(19,115,51));background-color:rgb(19,115,51);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(19,115,51))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.WFUiUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF13733300000000FF137333}.WFUiUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.WFUiUb .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF13733300000000FF137333}.WFUiUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.WFUiUb .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(19,115,51);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(19,115,51))}.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.WFUiUb .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(19,115,51);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(19,115,51))}.WFUiUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.WFUiUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.WFUiUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.WFUiUb .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.WFUiUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.WFUiUb .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(19,115,51)}.WFUiUb .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob:hover .VfPpkd-eHTEvd::before,.WFUiUb .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(19,115,51)}.WFUiUb .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(30,142,62)}.WFUiUb .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.WFUiUb .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(19,115,51)}.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(30,142,62)}.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(19,115,51)}.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(19,115,51)}.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(19,115,51)}.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(19,115,51)}.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(19,115,51)}.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.WFUiUb .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(19,115,51)}.WFUiUb .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#b1ddbd}.WFUiUb .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#b1ddbd}.WFUiUb .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#b1ddbd}.WFUiUb .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#b1ddbd}.WFUiUb .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(230,244,234)}.WFUiUb .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(19,115,51)}.WFUiUb .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(19,115,51)}.WFUiUb .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(19,115,51)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(30,142,62)}.WFUiUb .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.WFUiUb .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(30,142,62)}.WFUiUb .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.WFUiUb .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(30,142,62);background-color:var(--mdc-ripple-color,rgb(30,142,62))}.WFUiUb .U5B3me:not(:disabled){color:rgb(129,201,149)}.WFUiUb .U5B3me:not(:disabled):hover{color:rgb(129,201,149)}.WFUiUb .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.WFUiUb .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(129,201,149)}.WFUiUb .U5B3me .VfPpkd-Jh9lGc::before,.WFUiUb .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(129,201,149)}.WFUiUb .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(19,115,51)}.Mupove.bFjUmb-Ysl7Fe,.Mupove .bFjUmb-Ysl7Fe,.Mupove.CNpREd.bFjUmb-Ysl7Fe,.Mupove.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(243,232,253)}.Mupove.bFjUmb-Wvd9Cc,.Mupove .bFjUmb-Wvd9Cc,.Mupove.CNpREd.bFjUmb-Wvd9Cc,.Mupove.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(147,52,230)}.Mupove.bFjUmb-Tvm9db,.Mupove .bFjUmb-Tvm9db,.Mupove.CNpREd.bFjUmb-Tvm9db,.Mupove.CNpREd .bFjUmb-Tvm9db{background-color:rgb(118,39,187)}.Mupove.yxp05b-Wvd9Cc,.Mupove .yxp05b-Wvd9Cc,.Mupove.CNpREd.yxp05b-Wvd9Cc,.Mupove.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(147,52,230)}.Mupove.VnOHwf-Ysl7Fe,.Mupove .VnOHwf-Ysl7Fe,.Mupove.CNpREd.VnOHwf-Ysl7Fe,.Mupove.CNpREd .VnOHwf-Ysl7Fe{color:rgb(243,232,253);fill:rgb(243,232,253)}.Mupove.VnOHwf-Wvd9Cc,.Mupove .VnOHwf-Wvd9Cc,.Mupove.CNpREd.VnOHwf-Wvd9Cc,.Mupove.CNpREd .VnOHwf-Wvd9Cc{color:rgb(147,52,230);fill:rgb(147,52,230)}.Mupove.VnOHwf-Tvm9db,.Mupove .VnOHwf-Tvm9db,.Mupove.CNpREd.VnOHwf-Tvm9db,.Mupove.CNpREd .VnOHwf-Tvm9db{color:rgb(118,39,187);fill:rgb(118,39,187)}.Mupove.eL9Cfb,.Mupove .eL9Cfb,.Mupove.L5mE7d,.Mupove .L5mE7d,.Mupove.eL9Cfb:hover,.Mupove .eL9Cfb:hover,.Mupove.eL9Cfb:focus,.Mupove .eL9Cfb:focus,.Mupove.CNpREd.eL9Cfb,.Mupove.CNpREd .eL9Cfb,.Mupove.CNpREd.L5mE7d,.Mupove.CNpREd .L5mE7d,.Mupove.CNpREd.eL9Cfb:hover,.Mupove.CNpREd .eL9Cfb:hover,.Mupove.CNpREd.eL9Cfb:focus,.Mupove.CNpREd .eL9Cfb:focus{color:rgb(118,39,187)}.Mupove.L5mE7d:hover,.Mupove .L5mE7d:hover,.Mupove.L5mE7d:focus,.Mupove .L5mE7d:focus,.Mupove.L5mE7d:visited,.Mupove .L5mE7d:visited,.Mupove.CNpREd.L5mE7d:hover,.Mupove.CNpREd .L5mE7d:hover,.Mupove.CNpREd.L5mE7d:focus,.Mupove.CNpREd .L5mE7d:focus,.Mupove.CNpREd.L5mE7d:visited,.Mupove.CNpREd .L5mE7d:visited{color:rgb(147,52,230)}.Mupove .VUoKZ{background-color:rgb(243,232,253)}.Mupove .TRHLAc{background-color:rgb(147,52,230)}.Mupove .tgNIJf-Ysl7Fe:focus{border-color:rgb(243,232,253)}.Mupove .cjzpkc-Wvd9Cc:focus-within,.Mupove .tgNIJf-Wvd9Cc:focus{border-color:rgb(147,52,230)}.Mupove .u3bW4e .zZN2Lb-Wvd9Cc,.Mupove .zZN2Lb-Wvd9Cc:focus,.Mupove .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(147,52,230)}.Mupove .P3W0Dd-Ysl7Fe:focus,.Mupove.maXJsd:focus .P3W0Dd-Ysl7Fe,.Mupove .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(243,232,253)}.Mupove .VBEdtc-Wvd9Cc:hover,.Mupove.MymH0d:hover .VBEdtc-Wvd9Cc,.Mupove .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(147,52,230)}.Mupove.MymH0d:hover .UISY8d-Tvm9db,.Mupove.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.Mupove .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(147,52,230)}.Mupove .UISY8d-Ysl7Fe:hover,.Mupove.MymH0d:hover .UISY8d-Ysl7Fe,.Mupove .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(243,232,253)}.Mupove .mxmXhf{color:rgb(118,39,187);fill:rgb(118,39,187)}.Mupove .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.Mupove .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.Mupove .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.Mupove .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.Mupove .ZoT1D:focus-within.boxOzd,.Mupove .ZoT1D:focus-within.idtp4e,.Mupove .ZoT1D :focus-within.boxOzd,.Mupove .ZoT1D :focus-within.idtp4e{background-color:rgb(243,232,253)}.Mupove .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.Mupove .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.Mupove .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.Mupove .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.Mupove .ZoT1D:hover.j6KDAd,.Mupove .ZoT1D:hover.idtp4e,.Mupove .ZoT1D:hover .j6KDAd,.Mupove .ZoT1D:hover .idtp4e{background-color:rgb(243,232,253)}.Mupove .OGhwGf:hover,.Mupove .OGhwGf:focus{color:rgb(118,39,187)}.Mupove .ra2NV,.Mupove.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(147,52,230),transparent)}.Mupove .eumXzf:after{border-color:rgb(118,39,187)}.Mupove .zKHdkd .cXrdqd,.Mupove .kPBwDb{background-color:rgb(147,52,230)}.Mupove .zKHdkd .zHQkBf:not([disabled]):focus~.snByac,.Mupove .edhGSc.u3bW4e>.oJeWuf>.snByac{color:rgb(147,52,230)}.Mupove .bkIpNd .uHMk6b{border-color:rgb(243,232,253)}.Mupove .zJKIV .nQOrEb,.Mupove .zJKIV.RDPZE .nQOrEb,.Mupove .zJKIV.N2RpBe .Id5V1,.Mupove .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe .espmsb{border-color:rgb(147,52,230)}.Mupove .LsSwGf:not(.SWVgue):not(.RDPZE).N2RpBe>.MLPG7{border-color:rgb(147,52,230);opacity:.5}.Mupove .zJKIV.i9xfbb>.MbhUzd,.Mupove .zJKIV.u3bW4e>.MbhUzd,.Mupove .LsSwGf:not(.SWVgue).i9xfbb>.MbhUzd,.Mupove .LsSwGf:not(.SWVgue).u3bW4e>.MbhUzd{background-color:rgb(243,232,253)}.Mupove .HQ8yf:not(.RDPZE),.Mupove .HQ8yf:not(.RDPZE) a{color:rgb(147,52,230)}.Mupove .HQ8yf.u3bW4e .CeoRYc{background-color:rgba(147,52,230,.15)}.Mupove .HQ8yf .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(147,52,230,.25),rgba(147,52,230,.25) 80%,rgb(147,52,230) 100%)}.Mupove .uO32ac,.Mupove .ypv4re{border-bottom:1px solid rgb(147,52,230)}.Mupove .DqwBN:not(.RDPZE) .TpQm9d,.Mupove .l3F1ye:not(.RDPZE) .TpQm9d,.Mupove .YhQJj:not(.RDPZE) .TpQm9d,.Mupove .K2V86d:not(.RDPZE) .TpQm9d,.Mupove .An19kf:not(.RDPZE) .TpQm9d{color:rgb(118,39,187);fill:rgb(118,39,187)}.Mupove .DqwBN .TpQm9d,.Mupove .YhQJj .TpQm9d,.Mupove .K2V86d .TpQm9d,.Mupove .l3F1ye .TpQm9d,.Mupove .An19kf .TpQm9d{color:rgb(118,39,187);fill:rgb(118,39,187)}.Mupove .l3F1ye.j6PN2:not(.RDPZE) .TpQm9d{color:rgb(197,138,249);fill:rgb(197,138,249)}.Mupove .QkA63b:not(.RDPZE),.Mupove .Y5sE8d:not(.RDPZE){background-color:rgb(118,39,187)}.Mupove .An19kf:not(.RDPZE){background-color:rgb(243,232,253)}.Mupove .QkA63b:not(.RDPZE):hover,.Mupove .Y5sE8d:not(.RDPZE):hover,.Mupove .QkA63b:not(.RDPZE).u3bW4e,.Mupove .Y5sE8d:not(.RDPZE).u3bW4e{box-shadow:0 2px 1px -1px rgba(118,39,187,.2),0 1px 1px 0 rgba(118,39,187,.14),0 1px 3px 0 rgba(118,39,187,.12)}.Mupove .QkA63b:not(.RDPZE).iWO5td,.Mupove .Y5sE8d:not(.RDPZE).qs41qe{box-shadow:0 3px 5px -1px rgba(118,39,187,.2),0 6px 10px 0 rgba(118,39,187,.14),0 1px 18px 0 rgba(118,39,187,.12)}.Mupove .DqwBN:not(.RDPZE),.Mupove .YhQJj:not(.RDPZE),.Mupove .K2V86d:not(.RDPZE),.Mupove .l3F1ye:not(.RDPZE),.Mupove .An19kf:not(.RDPZE),.Mupove .BEAGS:not(.RDPZE),.Mupove .AeAAkf:not(.RDPZE){color:rgb(118,39,187)}.Mupove .l3F1ye.j6PN2:not(.RDPZE){color:rgb(197,138,249)}.Mupove .wwnMtb:not(.RDPZE),.Mupove .OZ6W0d:not(.RDPZE){color:rgb(118,39,187);fill:rgb(118,39,187)}.Mupove .wwnMtb:not(.RDPZE):hover,.Mupove .OZ6W0d:not(.RDPZE):hover{background-color:rgba(118,39,187,.08)}.Mupove .wwnMtb:not(.RDPZE).u3bW4e,.Mupove .OZ6W0d:not(.RDPZE).u3bW4e{background-color:rgba(118,39,187,.12)}.Mupove .wwnMtb:not(.RDPZE).u3bW4e:hover,.Mupove .OZ6W0d:not(.RDPZE).u3bW4e:hover{background-color:rgba(118,39,187,.16)}.Mupove .BEAGS.iWO5td,.Mupove .AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(118,39,187,.2),0 1px 1px 0 rgba(118,39,187,.14),0 1px 3px 0 rgba(118,39,187,.12)}.Mupove .DqwBN .MbhUzd,.Mupove .YhQJj .MbhUzd,.Mupove .K2V86d .MbhUzd,.Mupove .l3F1ye .MbhUzd,.Mupove .BEAGS .MbhUzd,.Mupove .AeAAkf .MbhUzd,.Mupove .An19kf .MbhUzd,.Mupove .OZ6W0d .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(118,39,187,.16),rgba(118,39,187,.16) 80%,rgba(118,39,187,0) 100%)}.Mupove .l3F1ye.j6PN2 .MbhUzd{background-image:radial-gradient(circle farthest-side,rgba(197,138,249,.16),rgba(197,138,249,.16) 80%,rgba(197,138,249,0) 100%)}.Mupove .AeAAkf:not(.RDPZE) .CeoRYc,.Mupove .BEAGS:not(.RDPZE) .CeoRYc,.Mupove .An19kf:not(.RDPZE) .CeoRYc,.Mupove .l3F1ye:not(.RDPZE) .CeoRYc,.Mupove .YhQJj:not(.RDPZE) .CeoRYc,.Mupove .K2V86d:not(.RDPZE) .CeoRYc,.Mupove .DqwBN:not(.RDPZE) .CeoRYc{background-color:rgb(118,39,187)}.Mupove .l3F1ye.j6PN2:not(.RDPZE) .CeoRYc{background-color:rgb(197,138,249)}.Mupove .AeAAkf:not(.RDPZE):hover,.Mupove .AeAAkf:not(.RDPZE).u3bW4e,.Mupove .BEAGS:not(.RDPZE):hover,.Mupove .BEAGS:not(.RDPZE).u3bW4e{border-color:rgba(147,52,230,.2)}.Mupove .DqwBN:not(.RDPZE):hover .CeoRYc,.Mupove .DqwBN:not(.RDPZE).u3bW4e .CeoRYc,.Mupove .YhQJj:not(.RDPZE):hover .CeoRYc,.Mupove .YhQJj:not(.RDPZE).u3bW4e .CeoRYc,.Mupove .K2V86d:not(.RDPZE):hover .CeoRYc,.Mupove .K2V86d:not(.RDPZE).u3bW4e .CeoRYc,.Mupove .An19kf:not(.RDPZE).u3bW4e .CeoRYc,.Mupove .l3F1ye:not(.RDPZE):hover .CeoRYc,.Mupove .l3F1ye:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(147,52,230)}.Mupove .l3F1ye.j6PN2:not(.RDPZE):hover .CeoRYc,.Mupove .l3F1ye.j6PN2:not(.RDPZE).u3bW4e .CeoRYc{background-color:rgb(197,138,249)}.Mupove .aiSeRd:not(.RDPZE).N2RpBe,.Mupove .aiSeRd:not(.RDPZE).B6Vhqe{border-color:rgb(147,52,230)}.Mupove .aiSeRd:not(.RDPZE):hover .MbhUzd,.Mupove .aiSeRd:not(.RDPZE):focus .MbhUzd,.Mupove .aiSeRd:not(.RDPZE).N2RpBe .MbhUzd,.Mupove .aiSeRd:not(.RDPZE).i9xfbb .MbhUzd{background-color:rgba(118,39,187,.08)}.Mupove .d7L4fc:hover .hYsg7c,.Mupove .NtlN8c:hover .hYsg7c{border-color:rgb(243,232,253)}.Mupove .d7L4fc:hover .MbhUzd,.Mupove .NtlN8c:hover .MbhUzd{background-color:rgba(118,39,187,.04)}.Mupove .d7L4fc .hYsg7c .nQOrEb,.Mupove .d7L4fc .hYsg7c.RDPZE .nQOrEb,.Mupove .d7L4fc .hYsg7c.N2RpBe .Id5V1{border-color:rgb(147,52,230)}.Mupove .d7L4fc .hYsg7c:not(.RDPZE).i9xfbb>.MbhUzd,.Mupove .d7L4fc .hYsg7c:not(.RDPZE).u3bW4e>.MbhUzd{background-color:rgba(118,39,187,.08)}.Mupove .SWVgue:not(.RDPZE).N2RpBe .espmsb{border-color:rgb(147,52,230)}.Mupove .SWVgue.RDPZE.N2RpBe .espmsb{border-color:#aa60eb}.Mupove .SWVgue:not(.RDPZE).N2RpBe .MLPG7{border-color:rgba(147,52,230,.3)}.Mupove .SWVgue.RDPZE.N2RpBe .MLPG7{border-color:#dbbbf7}.Mupove .SWVgue:not(.RDPZE).N2RpBe:hover .MbhUzd{background-color:rgba(147,52,230,.04)}.Mupove .SWVgue:not(.RDPZE).qs41qe .MbhUzd,.Mupove .SWVgue:not(.RDPZE).N2RpBe.u3bW4e .MbhUzd,.Mupove .SWVgue:not(.RDPZE).N2RpBe:focus .MbhUzd{background-color:rgba(147,52,230,.12)}.Mupove .HyS0Qd:not(.RDPZE) .zHQkBf,.Mupove .fWf7qe:not(.RDPZE) .tL9Q4c,.Mupove .D3oBEe:not(.RDPZE) .zHQkBf,.Mupove .AkVYk:not(.RDPZE) .tL9Q4c{caret-color:rgb(147,52,230)}.Mupove .HyS0Qd:not(.RDPZE) .cXrdqd,.Mupove .fWf7qe:not(.RDPZE) .cXrdqd,.Mupove .vnnr5e:not(.RDPZE) .cXrdqd{background-color:rgb(147,52,230)}.Mupove .D3oBEe:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before,.Mupove .AkVYk:not(.RDPZE).u3bW4e:not(.IYewr) .oJeWuf:before{border-color:rgb(147,52,230)}.Mupove .HyS0Qd:not(.RDPZE).u3bW4e .snByac,.Mupove .HyS0Qd input:not([disabled]):focus~.snByac,.Mupove .fWf7qe:not(.RDPZE).u3bW4e .snByac,.Mupove .D3oBEe:not(.RDPZE).u3bW4e .snByac,.Mupove .D3oBEe input:not([disabled]):focus~.snByac,.Mupove .AkVYk:not(.RDPZE).u3bW4e .snByac,.Mupove .vnnr5e:not(.RDPZE).u3bW4e .snByac{color:rgb(118,39,187)}.Mupove .ybOdnf:not(.RDPZE).iWO5td,.Mupove .ybOdnf:not(.RDPZE) .OA0qNb .LMgvRb[aria-selected=true],.Mupove .NqFm6:not(.RDPZE) .tWfTvb [role=option][aria-selected=true]{background-color:rgb(243,232,253)}.Mupove .RpYYWb:not(.RDPZE).fy1E5c .Ce1Y1c{color:rgb(147,52,230);fill:rgb(147,52,230)}.Mupove .mRipsb{background-color:rgb(147,52,230)}.Mupove .bJuVn.KKjvXb{background-color:rgb(118,39,187)}.Mupove .bJuVn.KKjvXb:before{background:linear-gradient(to top,rgb(118,39,187),transparent)}.Mupove .bJuVn.KKjvXb:after{background:linear-gradient(to bottom,rgb(118,39,187),transparent)}.Mupove .bJuVn.u3bW4e.KKjvXb.KKjvXb,.Mupove .bJuVn.KKjvXb.KKjvXb:hover{background-color:#7d29c7}.Mupove .bJuVn.u3bW4e.KKjvXb.KKjvXb:before,.Mupove .bJuVn.KKjvXb.KKjvXb:hover:before{background:linear-gradient(to top,#7d29c7,transparent)}.Mupove .bJuVn.u3bW4e.KKjvXb.KKjvXb:after,.Mupove .bJuVn.KKjvXb.KKjvXb:hover:after{background:linear-gradient(to bottom,#7d29c7,transparent)}.Mupove .pAlOFe{color:rgb(118,39,187);fill:rgb(118,39,187)}.Mupove .bDxw8b:not(:disabled){background-color:rgb(118,39,187)}.Mupove .FL3Khc:not(:disabled){color:rgb(118,39,187)}.Mupove .FL3Khc:not(:disabled):hover{color:rgb(118,39,187)}.Mupove .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Mupove .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(118,39,187)}.Mupove .FL3Khc .VfPpkd-Jh9lGc::before,.Mupove .FL3Khc .VfPpkd-Jh9lGc::after{background-color:rgb(118,39,187)}.Mupove .FL3Khc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Mupove .FL3Khc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(118,39,187)}.Mupove .n42Gr:not(:disabled){color:rgb(118,39,187)}.Mupove .n42Gr:not(:disabled):hover{color:rgb(118,39,187)}.Mupove .n42Gr:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Mupove .n42Gr:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(118,39,187)}.Mupove .n42Gr .VfPpkd-Jh9lGc::before,.Mupove .n42Gr .VfPpkd-Jh9lGc::after{background-color:rgb(118,39,187)}.Mupove .J5y29e:not(:disabled){color:rgb(118,39,187)}.Mupove .J5y29e:not(:disabled):hover{color:rgb(118,39,187)}.Mupove .J5y29e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Mupove .J5y29e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(118,39,187)}.Mupove .J5y29e .VfPpkd-Jh9lGc::before,.Mupove .J5y29e .VfPpkd-Jh9lGc::after{background-color:rgb(118,39,187)}.Mupove .LgeCif{color:rgb(118,39,187)}.Mupove .LgeCif:disabled{color:rgba(60,64,67,.38)}.Mupove .LgeCif .VfPpkd-Bz112c-Jh9lGc::before,.Mupove .LgeCif .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(118,39,187)}.Mupove .wlZwYd:not(:disabled){background-color:rgb(243,232,253)}.Mupove .wlZwYd:not(:disabled){color:rgb(118,39,187)}.Mupove .wlZwYd:not(:disabled):hover{color:rgb(118,39,187)}.Mupove .wlZwYd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Mupove .wlZwYd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(118,39,187)}.Mupove .wlZwYd .VfPpkd-Jh9lGc::before,.Mupove .wlZwYd .VfPpkd-Jh9lGc::after{background-color:rgb(118,39,187)}.Mupove .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}.Mupove .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Mupove .YJLdAc .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Mupove .YJLdAc .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(147,52,230);border-color:var(--mdc-checkbox-selected-icon-color,rgb(147,52,230));background-color:rgb(147,52,230);background-color:var(--mdc-checkbox-selected-icon-color,rgb(147,52,230))}@keyframes mdc-checkbox-fade-in-background-FF5F6368FF9334E600000000FF9334E6{0%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}50%{border-color:rgb(147,52,230);border-color:var(--mdc-checkbox-selected-icon-color,rgb(147,52,230));background-color:rgb(147,52,230);background-color:var(--mdc-checkbox-selected-icon-color,rgb(147,52,230))}}@keyframes mdc-checkbox-fade-out-background-FF5F6368FF9334E600000000FF9334E6{0%,80%{border-color:rgb(147,52,230);border-color:var(--mdc-checkbox-selected-icon-color,rgb(147,52,230));background-color:rgb(147,52,230);background-color:var(--mdc-checkbox-selected-icon-color,rgb(147,52,230))}100%{border-color:rgb(95,99,104);border-color:var(--mdc-checkbox-unselected-icon-color,rgb(95,99,104));background-color:transparent}}.Mupove .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF5F6368FF9334E600000000FF9334E6}.Mupove .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF5F6368FF9334E600000000FF9334E6}.Mupove .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-hover-icon-color,rgb(32,33,36));background-color:transparent}.Mupove .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Mupove .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Mupove .YJLdAc:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(118,39,187);border-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(118,39,187));background-color:rgb(118,39,187);background-color:var(--mdc-checkbox-selected-hover-icon-color,rgb(118,39,187))}.Mupove .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF7627BB00000000FF7627BB}.Mupove .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF7627BB00000000FF7627BB}.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-focus-icon-color,rgb(32,33,36));background-color:transparent}.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(118,39,187);border-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(118,39,187));background-color:rgb(118,39,187);background-color:var(--mdc-checkbox-selected-focus-icon-color,rgb(118,39,187))}.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF7627BB00000000FF7627BB}.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF7627BB00000000FF7627BB}.Mupove .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}.Mupove .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:rgb(118,39,187);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(118,39,187));background-color:rgb(118,39,187);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(118,39,187))}@keyframes mdc-checkbox-fade-in-background-FF202124FF7627BB00000000FF7627BB{0%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}50%{border-color:rgb(118,39,187);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(118,39,187));background-color:rgb(118,39,187);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(118,39,187))}}@keyframes mdc-checkbox-fade-out-background-FF202124FF7627BB00000000FF7627BB{0%,80%{border-color:rgb(118,39,187);border-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(118,39,187));background-color:rgb(118,39,187);background-color:var(--mdc-checkbox-selected-pressed-icon-color,rgb(118,39,187))}100%{border-color:rgb(32,33,36);border-color:var(--mdc-checkbox-unselected-pressed-icon-color,rgb(32,33,36));background-color:transparent}}.Mupove .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-in-background-FF202124FF7627BB00000000FF7627BB}.Mupove .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.Mupove .YJLdAc:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{animation-name:mdc-checkbox-fade-out-background-FF202124FF7627BB00000000FF7627BB}.Mupove .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.Mupove .YJLdAc.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(118,39,187);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(118,39,187))}.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.Mupove .YJLdAc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:rgb(118,39,187);background-color:var(--mdc-checkbox-selected-hover-state-layer-color,rgb(118,39,187))}.Mupove .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.Mupove .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.Mupove .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.Mupove .sPi0ob.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::after,.Mupove .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before,.Mupove .sPi0ob:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::after{background-color:rgb(118,39,187)}.Mupove .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob:hover .VfPpkd-eHTEvd::before,.Mupove .sPi0ob:hover .VfPpkd-eHTEvd::after{background-color:rgb(118,39,187)}.Mupove .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob:not(:disabled):active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(147,52,230)}.Mupove .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::before,.Mupove .sPi0ob:not(:disabled):active .VfPpkd-eHTEvd::after{background-color:rgb(118,39,187)}.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(147,52,230)}.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(118,39,187)}.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(118,39,187)}.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(118,39,187)}.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(118,39,187)}.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(118,39,187)}.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.Mupove .dcwaj.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(118,39,187)}.Mupove .dcwaj:enabled .VfPpkd-l6JLsf::after{background:#cea2f7}.Mupove .dcwaj:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:#cea2f7}.Mupove .dcwaj:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:#cea2f7}.Mupove .dcwaj:enabled:active .VfPpkd-l6JLsf::after{background:#cea2f7}.Mupove .g0jqJf .VfPpkd-OkbHre.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(243,232,253)}.Mupove .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(118,39,187)}.Mupove .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(118,39,187)}.Mupove .g0jqJf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(118,39,187)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(147,52,230)}.Mupove .I2Xlzb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after,.Mupove .mCP2Kb .CFILmd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(147,52,230)}.Mupove .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::before,.Mupove .mCP2Kb .eJy6Bb .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(147,52,230);background-color:var(--mdc-ripple-color,rgb(147,52,230))}.Mupove .U5B3me:not(:disabled){color:rgb(197,138,249)}.Mupove .U5B3me:not(:disabled):hover{color:rgb(197,138,249)}.Mupove .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Mupove .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(197,138,249)}.Mupove .U5B3me .VfPpkd-Jh9lGc::before,.Mupove .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(197,138,249)}.Mupove .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(118,39,187)}.kYtXye.bFjUmb-Ysl7Fe,.kYtXye .bFjUmb-Ysl7Fe,.kYtXye.CNpREd.bFjUmb-Ysl7Fe,.kYtXye.CNpREd .bFjUmb-Ysl7Fe{background-color:rgb(232,240,254)}.kYtXye.bFjUmb-Wvd9Cc,.kYtXye .bFjUmb-Wvd9Cc,.kYtXye.CNpREd.bFjUmb-Wvd9Cc,.kYtXye.CNpREd .bFjUmb-Wvd9Cc{background-color:rgb(26,115,232)}.kYtXye.bFjUmb-Tvm9db,.kYtXye .bFjUmb-Tvm9db,.kYtXye.CNpREd.bFjUmb-Tvm9db,.kYtXye.CNpREd .bFjUmb-Tvm9db{background-color:rgb(24,90,188)}.kYtXye.yxp05b-Wvd9Cc,.kYtXye .yxp05b-Wvd9Cc,.kYtXye.CNpREd.yxp05b-Wvd9Cc,.kYtXye.CNpREd .yxp05b-Wvd9Cc{border-color:rgb(26,115,232)}.kYtXye.VnOHwf-Ysl7Fe,.kYtXye .VnOHwf-Ysl7Fe,.kYtXye.CNpREd.VnOHwf-Ysl7Fe,.kYtXye.CNpREd .VnOHwf-Ysl7Fe{color:rgb(232,240,254);fill:rgb(232,240,254)}.kYtXye.VnOHwf-Wvd9Cc,.kYtXye .VnOHwf-Wvd9Cc,.kYtXye.CNpREd.VnOHwf-Wvd9Cc,.kYtXye.CNpREd .VnOHwf-Wvd9Cc{color:rgb(26,115,232);fill:rgb(26,115,232)}.kYtXye.VnOHwf-Tvm9db,.kYtXye .VnOHwf-Tvm9db,.kYtXye.CNpREd.VnOHwf-Tvm9db,.kYtXye.CNpREd .VnOHwf-Tvm9db{color:rgb(24,90,188);fill:rgb(24,90,188)}.kYtXye.eL9Cfb,.kYtXye .eL9Cfb,.kYtXye.L5mE7d,.kYtXye .L5mE7d,.kYtXye.eL9Cfb:hover,.kYtXye .eL9Cfb:hover,.kYtXye.eL9Cfb:focus,.kYtXye .eL9Cfb:focus,.kYtXye.CNpREd.eL9Cfb,.kYtXye.CNpREd .eL9Cfb,.kYtXye.CNpREd.L5mE7d,.kYtXye.CNpREd .L5mE7d,.kYtXye.CNpREd.eL9Cfb:hover,.kYtXye.CNpREd .eL9Cfb:hover,.kYtXye.CNpREd.eL9Cfb:focus,.kYtXye.CNpREd .eL9Cfb:focus{color:rgb(24,90,188)}.kYtXye.L5mE7d:hover,.kYtXye .L5mE7d:hover,.kYtXye.L5mE7d:focus,.kYtXye .L5mE7d:focus,.kYtXye.L5mE7d:visited,.kYtXye .L5mE7d:visited,.kYtXye.CNpREd.L5mE7d:hover,.kYtXye.CNpREd .L5mE7d:hover,.kYtXye.CNpREd.L5mE7d:focus,.kYtXye.CNpREd .L5mE7d:focus,.kYtXye.CNpREd.L5mE7d:visited,.kYtXye.CNpREd .L5mE7d:visited{color:rgb(26,115,232)}.kYtXye .VUoKZ{background-color:rgb(232,240,254)}.kYtXye .TRHLAc{background-color:rgb(26,115,232)}.kYtXye .tgNIJf-Ysl7Fe:focus{border-color:rgb(232,240,254)}.kYtXye .cjzpkc-Wvd9Cc:focus-within,.kYtXye .tgNIJf-Wvd9Cc:focus{border-color:rgb(26,115,232)}.kYtXye .u3bW4e .zZN2Lb-Wvd9Cc,.kYtXye .zZN2Lb-Wvd9Cc:focus,.kYtXye .maXJsd:focus .zZN2Lb-Wvd9Cc{color:rgb(26,115,232)}.kYtXye .P3W0Dd-Ysl7Fe:focus,.kYtXye.maXJsd:focus .P3W0Dd-Ysl7Fe,.kYtXye .maXJsd:focus .P3W0Dd-Ysl7Fe{background-color:rgb(232,240,254)}.kYtXye .VBEdtc-Wvd9Cc:hover,.kYtXye.MymH0d:hover .VBEdtc-Wvd9Cc,.kYtXye .MymH0d:hover .VBEdtc-Wvd9Cc{color:rgb(26,115,232)}.kYtXye.MymH0d:hover .UISY8d-Tvm9db,.kYtXye.CNpREd.MymH0d:hover .UISY8d-Tvm9db,.kYtXye .MymH0d:hover .UISY8d-Tvm9db{background-color:rgb(26,115,232)}.kYtXye .UISY8d-Ysl7Fe:hover,.kYtXye.MymH0d:hover .UISY8d-Ysl7Fe,.kYtXye .MymH0d:hover .UISY8d-Ysl7Fe{background-color:rgb(232,240,254)}.kYtXye .mxmXhf{color:rgb(24,90,188);fill:rgb(24,90,188)}.kYtXye .tUJKGd:not(.xp2dJ):focus-within.boxOzd,.kYtXye .tUJKGd:not(.xp2dJ):focus-within.idtp4e,.kYtXye .tUJKGd:not(.xp2dJ) :focus-within.boxOzd,.kYtXye .tUJKGd:not(.xp2dJ) :focus-within.idtp4e,.kYtXye .ZoT1D:focus-within.boxOzd,.kYtXye .ZoT1D:focus-within.idtp4e,.kYtXye .ZoT1D :focus-within.boxOzd,.kYtXye .ZoT1D :focus-within.idtp4e{background-color:rgb(232,240,254)}.kYtXye .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.j6KDAd,.kYtXye .tUJKGd:not(.xp2dJ):not(.rZXyy):hover.idtp4e,.kYtXye .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .j6KDAd,.kYtXye .tUJKGd:not(.xp2dJ):not(.rZXyy):hover .idtp4e,.kYtXye .ZoT1D:hover.j6KDAd,.kYtXye .ZoT1D:hover.idtp4e,.kYtXye .ZoT1D:hover .j6KDAd,.kYtXye .ZoT1D:hover .idtp4e{background-color:rgb(232,240,254)}.kYtXye .OGhwGf:hover,.kYtXye .OGhwGf:focus{color:rgb(24,90,188)}.kYtXye .ra2NV,.kYtXye.ra2NV.ra2NV{background-image:radial-gradient(25rem 18.75rem ellipse at bottom right,rgb(26,115,232),transparent)}.kYtXye .eumXzf:after{border-color:rgb(24,90,188)}.kYtXye .uO32ac,.kYtXye .ypv4re{border-bottom:1px solid rgb(26,115,232)}.kYtXye .U5B3me:not(:disabled){color:rgb(138,180,248)}.kYtXye .U5B3me:not(:disabled):hover{color:rgb(138,180,248)}.kYtXye .U5B3me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.kYtXye .U5B3me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(138,180,248)}.kYtXye .U5B3me .VfPpkd-Jh9lGc::before,.kYtXye .U5B3me .VfPpkd-Jh9lGc::after{background-color:rgb(138,180,248)}.kYtXye .AzAT4d .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(24,90,188)}html{height:100%}body{height:100%;-moz-osx-font-smoothing:grayscale;color:rgba(0,0,0,.87);font-family:Roboto,RobotoDraft,Helvetica,Arial,sans-serif;margin:0;-moz-text-size-adjust:100%;-moz-text-size-adjust:100%;text-size-adjust:100%}textarea{font-family:Roboto,RobotoDraft,Helvetica,Arial,sans-serif}a{text-decoration:none;color:#2962ff}img{border:none}#apps-debug-tracers{display:none}html{overflow:visible}body{overflow:visible;overflow-y:scroll}@keyframes quantumWizBoxInkSpread{0%{transform:translate(-50%,-50%) scale(0.2)}to{transform:translate(-50%,-50%) scale(2.2)}}@keyframes quantumWizIconFocusPulse{0%{transform:translate(-50%,-50%) scale(1.5);opacity:0}to{transform:translate(-50%,-50%) scale(2);opacity:1}}@keyframes quantumWizRadialInkSpread{0%{transform:scale(1.5);opacity:0}to{transform:scale(2.5);opacity:1}}@keyframes quantumWizRadialInkFocusPulse{0%{transform:scale(2);opacity:0}to{transform:scale(2.5);opacity:1}}.mUbCce{-moz-user-select:none;-moz-transition:background .3s;transition:background .3s;border:0;-moz-border-radius:50%;border-radius:50%;cursor:pointer;display:inline-block;flex-shrink:0;height:48px;outline:none;overflow:hidden;position:relative;text-align:center;width:48px;z-index:0}.mUbCce>.TpQm9d{height:48px;width:48px}.YYBxpf{-moz-border-radius:0;border-radius:0;overflow:visible}.fKz7Od{color:rgba(0,0,0,.54);fill:rgba(0,0,0,.54)}.p9Nwte{color:rgba(255,255,255,.75);fill:rgba(255,255,255,.75)}.fKz7Od.u3bW4e{background-color:rgba(0,0,0,.12)}.p9Nwte.u3bW4e{background-color:rgba(204,204,204,.25)}.YYBxpf.u3bW4e{background-color:transparent}.VTBa7b{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s,-webkit-transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,-webkit-transform 0s ease .2s;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.YYBxpf.u3bW4e .VTBa7b{-moz-animation:quantumWizIconFocusPulse .7s infinite alternate;animation:quantumWizIconFocusPulse .7s infinite alternate;height:100%;left:50%;top:50%;width:100%;visibility:visible}.mUbCce.qs41qe .VTBa7b{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.mUbCce.qs41qe.M9Bg4d .VTBa7b{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1);transition:opacity .2s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1)}.mUbCce.j7nIZb .VTBa7b{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);visibility:visible}.fKz7Od .VTBa7b{background-image:radial-gradient(circle farthest-side,rgba(0,0,0,.12),rgba(0,0,0,.12) 80%,rgba(0,0,0,0) 100%)}.p9Nwte .VTBa7b{background-image:radial-gradient(circle farthest-side,rgba(204,204,204,.25),rgba(204,204,204,.25) 80%,rgba(204,204,204,0) 100%)}.mUbCce.RDPZE{color:rgba(0,0,0,.26);fill:rgba(0,0,0,.26);cursor:default}.p9Nwte.RDPZE{color:rgba(255,255,255,0.502);fill:rgba(255,255,255,0.502)}.xjKiLb{position:relative;top:50%}.xjKiLb>span{display:inline-block;position:relative}.ettIx{width:300px}.cnOaDb{overflow-wrap:break-word;position:relative}.cnOaDb.vTcY1d{padding-top:24px}.cnOaDb.sgOJyf{padding-bottom:24px}.T2Ybvb{outline:none}.T2Ybvb:empty:before{content:"\0000a0"}.nZC2Ae,.iSSROb{color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;left:0;pointer-events:none;position:absolute;right:0}.cnOaDb.vTcY1d .nZC2Ae{top:24px}.cnOaDb.sgOJyf .nZC2Ae{bottom:24px}.iSSROb{top:0}.nZC2Ae{transform-origin:bottom left;transition-property:color,-webkit-transform;transition-property:color,transform;transition-property:color,transform,-webkit-transform;transition:all .3s cubic-bezier(0.4,0,0.2,1)}.ettIx.u3bW4e:not(.RDPZE) .nZC2Ae{color:#4285f4}.ettIx.u3bW4e:not(.RDPZE) .nZC2Ae,.ettIx.CDELXb .nZC2Ae{transform:scale(0.75) translateY(-39px)}.ettIx.u3bW4e:not(.RDPZE) .cnOaDb.sgOJyf .nZC2Ae,.ettIx.CDELXb .cnOaDb.sgOJyf .nZC2Ae{transform:scale(0.75) translateY(39px)}.ettIx.CDELXb .iSSROb{display:none}.ettIx.RDPZE .T2Ybvb,.ettIx.RDPZE .nZC2Ae,.ettIx.RDPZE .iSSROb{opacity:.54}.tsIGMc,.PfAg4{bottom:-2px;left:0;margin:0;padding:0;position:absolute;width:100%}.cnOaDb.sgOJyf .tsIGMc,.cnOaDb.sgOJyf .PfAg4{bottom:22px}.tsIGMc{background-color:rgba(0,0,0,.12);height:1px}.ettIx.RDPZE .tsIGMc{background:none;border-bottom:1px dotted rgba(0,0,0,.12)}.PfAg4{animation:RemoveUnderline .3s cubic-bezier(0.4,0,0.2,1);background-color:#4285f4;height:2px;transform:scaleX(0)}@keyframes RemoveUnderline{0%{opacity:1;-moz-transform:scaleX(1);transform:scaleX(1)}to{opacity:0;-moz-transform:scaleX(1);transform:scaleX(1)}}.ettIx.u3bW4e:not(.RDPZE) .PfAg4{animation:AddUnderline .3s cubic-bezier(0.4,0,0.2,1);transform:scaleX(1)}@keyframes AddUnderline{0%{-moz-transform:scaleX(0);transform:scaleX(0)}to{-moz-transform:scaleX(1);transform:scaleX(1)}}.qmMNRc{color:rgba(0,0,0,.54);height:34px;margin-top:2px;width:36px}.Erb9le:not(.RDPZE) .qmMNRc:hover,.Erb9le:not(.RDPZE) .qmMNRc.y7OZL{color:rgba(0,0,0,.87)}.Erb9le:not(.RDPZE) .qmMNRc.y7OZL{background-color:#e0e0e0;-moz-border-radius:2px;border-radius:2px}.FKF6mc,.FKF6mc:focus{display:block;outline:none;text-decoration:none}.FKF6mc:visited{fill:inherit;stroke:inherit}.U26fgb.u3bW4e{outline:1px solid transparent}.DPvwYc{font-family:"Material Icons Extended";font-weight:normal;font-style:normal;font-size:24px;line-height:1;letter-spacing:normal;text-rendering:optimizeLegibility;text-transform:none;display:inline-block;word-wrap:normal;direction:ltr;font-feature-settings:"liga" 1}html[dir="rtl"] .sm8sCf{-moz-transform:scaleX(-1);transform:scaleX(-1);filter:FlipH}.UQuaGc{transition:box-shadow 280ms cubic-bezier(0.4,0,0.2,1);-moz-user-select:none;-moz-transition:background .2s .1s;transition:background .2s .1s;border:0;-moz-border-radius:4px;border-radius:4px;color:#5f6368;cursor:pointer;display:inline-block;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:14px;font-weight:500;letter-spacing:.25px;line-height:36px;text-decoration:none;text-transform:none;min-width:auto;outline:none;overflow:hidden;position:relative;text-align:center;z-index:0}.UQuaGc.qs41qe{transition:box-shadow 280ms cubic-bezier(0.4,0,0.2,1)}.DRsGyd{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:13px;font-weight:500;letter-spacing:.25px;line-height:24px;text-decoration:none;text-transform:none}.UQuaGc.TuHiFd{width:100%}.TuHiFd .l4V7wb{justify-content:center}.Y5sE8d{background:#1a73e8;color:#fff}.UQuaGc.Y5sE8d.qs41qe{box-shadow:0 3px 5px -1px rgba(26,115,232,0.2),0 6px 10px 0 rgba(26,115,232,0.141),0 1px 18px 0 rgba(26,115,232,0.122)}.An19kf{background:#e8f0fe;color:#1967d2}.UQuaGc.An19kf.qs41qe{box-shadow:0 3px 5px -1px rgba(0,0,0,0.2),0 6px 10px 0 rgba(0,0,0,0.141),0 1px 18px 0 rgba(0,0,0,0.122)}.l3F1ye,.l3F1ye .TpQm9d{color:#1a73e8}.j6PN2,.j6PN2 .TpQm9d{color:#e8eaed}.j6PN2.l3F1ye,.j6PN2.l3F1ye .TpQm9d{color:#8ab4f8}.j6PN2.l3F1ye.qs41qe,.j6PN2.l3F1ye.qs41qe .TpQm9d{color:#aecbfa}.AeAAkf{border:1px #dadce0 solid;box-sizing:border-box;color:#1a73e8;height:36px;line-height:34px}.AeAAkf.DRsGyd{height:24px;line-height:22px}.YWP0Id.UQuaGc{align-items:center;box-sizing:border-box;display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;height:auto;line-height:normal;min-height:36px}.YWP0Id.DRsGyd{min-height:24px}.AeAAkf.qs41qe{box-shadow:0 2px 1px -1px rgba(26,115,232,0.2),0 1px 1px 0 rgba(26,115,232,0.141),0 1px 3px 0 rgba(26,115,232,0.122);border:none}.Y5sE8d .TpQm9d,.Y5sE8d .TpQm9d:hover,.Y5sE8d .TpQm9d:link,.Y5sE8d .TpQm9d:visited{color:#fff}.An19kf .TpQm9d,.An19kf .TpQm9d:hover,.An19kf .TpQm9d:link,.An19kf .TpQm9d:visited{color:#1967d2}.YhQJj{box-shadow:0 2px 1px -1px rgba(0,0,0,0.2),0 1px 1px 0 rgba(0,0,0,0.141),0 1px 3px 0 rgba(0,0,0,0.122);background-color:#fff;color:#1a73e8}.YhQJj.qs41qe{box-shadow:0 3px 5px -1px rgba(0,0,0,0.2),0 6px 10px 0 rgba(0,0,0,0.141),0 1px 18px 0 rgba(0,0,0,0.122)}.e19J0b{position:absolute;top:0;right:0;bottom:0;left:0;background-color:#5f6368;opacity:0}.j6PN2 .e19J0b{background-color:#e8eaed}.j6PN2.l3F1ye .e19J0b{background-color:#8ab4f8}.Y5sE8d .e19J0b{background-color:#fff}.An19kf .e19J0b{background-color:#1a73e8}.l3F1ye .e19J0b,.AeAAkf .e19J0b,.YhQJj .e19J0b{background-color:#4285f4}.UQuaGc:hover .e19J0b{opacity:0.04}.AeAAkf:hover{border-color:#d2e3fc}.Y5sE8d:hover{box-shadow:0 2px 1px -1px rgba(26,115,232,0.2),0 1px 1px 0 rgba(26,115,232,0.141),0 1px 3px 0 rgba(26,115,232,0.122)}.An19kf:hover{box-shadow:0 2px 1px -1px rgba(0,0,0,0.2),0 1px 1px 0 rgba(0,0,0,0.141),0 1px 3px 0 rgba(0,0,0,0.122)}.j6PN2:hover .e19J0b{opacity:0.04}.Y5sE8d:hover .e19J0b{opacity:0.08}.UQuaGc.u3bW4e .e19J0b{opacity:0.12}.l3F1ye.u3bW4e,.l3F1ye.u3bW4e .TpQm9d{color:#1967d2}.j6PN2.l3F1ye.u3bW4e,.j6PN2.l3F1ye.u3bW4e .TpQm9d{color:#8ab4f8}.j6PN2.u3bW4e .e19J0b{opacity:0.12}.An19kf.u3bW4e,.An19kf.u3bW4e .TpQm9d,.An19kf.u3bW4e .TpQm9d:hover,.An19kf.u3bW4e .TpQm9d:link,.An19kf.u3bW4e .TpQm9d:visited{color:#185abc}.AeAAkf.u3bW4e{color:#1967d2;border-color:#d2e3fc}.YhQJj.u3bW4e{color:#1967d2}.Y5sE8d.u3bW4e .e19J0b{opacity:0.24}.UQuaGc.u3bW4e:hover .e19J0b{opacity:0.155}.j6PN2.u3bW4e:hover .e19J0b{opacity:0.155}.Y5sE8d.u3bW4e:hover .e19J0b{opacity:0.3}.UQuaGc.RDPZE .e19J0b{opacity:0}.Fvio9d{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,-webkit-transform 0s ease .2s;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.UQuaGc.qs41qe .Fvio9d{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.UQuaGc.qs41qe.M9Bg4d .Fvio9d{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1)}.UQuaGc.j7nIZb .Fvio9d{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);visibility:visible}.kCyAyd .Fvio9d{background-image:radial-gradient(circle farthest-side,rgba(0,0,0,.12),rgba(0,0,0,.12) 80%,rgba(0,0,0,0) 100%)}.l3F1ye .Fvio9d,.AeAAkf .Fvio9d,.YhQJj .Fvio9d{background-image:radial-gradient(circle farthest-side,rgba(66,133,244,0.161),rgba(66,133,244,0.161) 80%,rgba(66,133,244,0) 100%)}.An19kf .Fvio9d{background-image:radial-gradient(circle farthest-side,rgba(26,115,232,0.161),rgba(26,115,232,0.161) 80%,rgba(26,115,232,0) 100%)}.j6PN2 .Fvio9d{background-image:radial-gradient(circle farthest-side,rgba(232,234,237,0.161),rgba(232,234,237,0.161) 80%,rgba(232,234,237,0) 100%)}.j6PN2.l3F1ye .Fvio9d{background-image:radial-gradient(circle farthest-side,rgba(174,203,250,0.161),rgba(174,203,250,0.161) 80%,rgba(174,203,250,0) 100%)}.Y5sE8d .Fvio9d{background-image:radial-gradient(circle farthest-side,rgba(255,255,255,0.322),rgba(255,255,255,0.322) 80%,rgba(255,255,255,0) 100%)}.UQuaGc.RDPZE{-moz-box-shadow:none;box-shadow:none;color:rgba(0,0,0,.38);cursor:default;fill:rgba(0,0,0,.38)}.j6PN2.RDPZE{color:rgba(255,255,255,.38);fill:rgba(255,255,255,.38)}.AeAAkf.RDPZE,.AeAAkf.RDPZE:hover{border-color:rgba(0,0,0,.12)}.Y5sE8d.RDPZE,.YhQJj.RDPZE,.An19kf.RDPZE{background:rgba(0,0,0,.12)}.l4V7wb{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;position:relative}.l4V7wb .NPEfkd{display:inline-block;margin:0}.kCyAyd .l4V7wb,.l3F1ye .l4V7wb{padding:0 8px}.AeAAkf .l4V7wb{padding:0 23px}.AeAAkf.qs41qe .l4V7wb{padding:1px 24px}.Y5sE8d .l4V7wb,.YhQJj .l4V7wb,.An19kf .l4V7wb{padding:0 24px}.DRsGyd.AeAAkf .l4V7wb{padding:0 11px}.DRsGyd.AeAAkf.qs41qe .l4V7wb{padding:1px 12px}.DRsGyd.Y5sE8d .l4V7wb,.DRsGyd.YhQJj .l4V7wb{padding:0 12px}.l4V7wb.cd29Sd{padding:0 16px 0 12px}.l4V7wb.cd29Sd.olttVd{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-orient:horizontal;box-orient:horizontal;flex-direction:row-reverse;padding:0 12px 0 16px}.AeAAkf.qs41qe .cd29Sd.l4V7wb{padding:1px 16px 1px 12px}.AeAAkf.qs41qe .cd29Sd.olttVd.l4V7wb{padding:1px 12px 1px 16px}.AeAAkf .cd29Sd.l4V7wb{padding:0 15px 0 11px}.AeAAkf .cd29Sd.olttVd.l4V7wb{padding:0 0;padding:0 -moz-calc(12px - 1px) 0 -moz-calc(16px - 1px);padding:0 calc(12px - 1px) 0 calc(16px - 1px)}.E6FpNe{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;color:currentcolor;fill:currentcolor;margin-right:8px}.l4V7wb.olttVd .E6FpNe{margin-left:8px;margin-right:0}.Y5FYJe{-moz-user-select:none;-moz-transition:background .3s;transition:background .3s;border:0;-moz-border-radius:50%;border-radius:50%;cursor:pointer;display:inline-block;flex-shrink:0;height:48px;outline:none;overflow:hidden;position:relative;text-align:center;width:48px;z-index:0}.Y5FYJe>.TpQm9d{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:48px;width:48px}.L23pJb{overflow:visible}.Y5FYJe:hover{background-color:rgba(95,99,104,0.039)}.Y5FYJe.RDPZE:hover{background-color:transparent}.VsxsTb:hover{background-color:rgba(232,234,237,0.039)}.OZ6W0d:hover{background-color:rgba(66,133,244,0.039)}.cjq2Db{color:#5f6368;fill:#5f6368}.VsxsTb{color:#e8eaed;fill:#e8eaed}.OZ6W0d{color:#1a73e8;fill:#1a73e8}.cjq2Db.u3bW4e{background-color:rgba(95,99,104,0.122)}.cjq2Db.u3bW4e:hover{background-color:rgba(95,99,104,0.157)}.VsxsTb.u3bW4e{background-color:rgba(232,234,237,0.122)}.VsxsTb.u3bW4e:hover{background-color:rgba(232,234,237,0.157)}.OZ6W0d.u3bW4e{background-color:rgba(66,133,244,0.122)}.OZ6W0d.u3bW4e:hover{background-color:rgba(66,133,244,0.157)}.L23pJb.u3bW4e{background-color:transparent}.PDXc1b{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,-webkit-transform 0s ease .2s;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.L23pJb.u3bW4e .PDXc1b{-moz-animation:quantumWizIconFocusPulse .7s infinite alternate;animation:quantumWizIconFocusPulse .7s infinite alternate;height:100%;left:50%;top:50%;width:100%;visibility:visible}.Y5FYJe.qs41qe .PDXc1b{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.Y5FYJe.qs41qe.M9Bg4d .PDXc1b{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1)}.Y5FYJe.j7nIZb .PDXc1b{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);visibility:visible}.cjq2Db .PDXc1b{background-image:radial-gradient(circle farthest-side,rgba(95,99,104,0.161),rgba(95,99,104,0.161) 80%,rgba(95,99,104,0) 100%)}.VsxsTb .PDXc1b{background-image:radial-gradient(circle farthest-side,rgba(255,255,255,0.161),rgba(255,255,255,0.161) 80%,rgba(255,255,255,0) 100%)}.OZ6W0d .PDXc1b{background-image:radial-gradient(circle farthest-side,rgba(66,133,244,0.161),rgba(66,133,244,0.161) 80%,rgba(66,133,244,0) 100%)}.Y5FYJe.RDPZE{color:#9aa0a6;fill:#9aa0a6;cursor:default}.VsxsTb.RDPZE{color:rgba(255,255,255,.38);fill:rgba(255,255,255,.38)}.XuQwKc{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:100%;justify-content:center;position:relative;width:100%}.GmuOkf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;position:relative}.O0WRkf{-moz-user-select:none;-moz-transition:background .2s .1s;transition:background .2s .1s;border:0;-moz-border-radius:3px;border-radius:3px;cursor:pointer;display:inline-block;font-size:14px;font-weight:500;min-width:4em;outline:none;overflow:hidden;position:relative;text-align:center;text-transform:uppercase;z-index:0}.A9jyad{font-size:13px;line-height:16px}.zZhnYe{-moz-transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);background:#dfdfdf;-moz-box-shadow:0px 2px 2px 0px rgba(0,0,0,.14),0px 3px 1px -2px rgba(0,0,0,.12),0px 1px 5px 0px rgba(0,0,0,.2);box-shadow:0px 2px 2px 0px rgba(0,0,0,.14),0px 3px 1px -2px rgba(0,0,0,.12),0px 1px 5px 0px rgba(0,0,0,.2)}.zZhnYe.qs41qe{-moz-transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);-moz-transition:background .8s;transition:background .8s;-moz-box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2)}.e3Duub,.e3Duub a,.e3Duub a:hover,.e3Duub a:link,.e3Duub a:visited{background:#4285f4;color:#fff}.HQ8yf,.HQ8yf a{color:#4285f4}.UxubU,.UxubU a{color:#fff}.ZFr60d{position:absolute;top:0;right:0;bottom:0;left:0;background-color:transparent}.O0WRkf.u3bW4e .ZFr60d{background-color:rgba(0,0,0,.12)}.UxubU.u3bW4e .ZFr60d{background-color:rgba(255,255,255,.3)}.e3Duub.u3bW4e .ZFr60d{background-color:rgba(0,0,0,0.122)}.HQ8yf.u3bW4e .ZFr60d{background-color:rgba(66,133,244,.15)}.Vwe4Vb{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s,-webkit-transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,-webkit-transform 0s ease .2s;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.O0WRkf.qs41qe .Vwe4Vb{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.O0WRkf.qs41qe.M9Bg4d .Vwe4Vb{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1);transition:opacity .2s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1)}.O0WRkf.j7nIZb .Vwe4Vb{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);visibility:visible}.oG5Srb .Vwe4Vb,.zZhnYe .Vwe4Vb{background-image:radial-gradient(circle farthest-side,rgba(0,0,0,.12),rgba(0,0,0,.12) 80%,rgba(0,0,0,0) 100%)}.HQ8yf .Vwe4Vb{background-image:radial-gradient(circle farthest-side,rgba(66,133,244,.25),rgba(66,133,244,.25) 80%,rgba(66,133,244,0) 100%)}.e3Duub .Vwe4Vb{background-image:radial-gradient(circle farthest-side,#3367d6,#3367d6 80%,rgba(51,103,214,0) 100%)}.UxubU .Vwe4Vb{background-image:radial-gradient(circle farthest-side,rgba(255,255,255,.3),rgba(255,255,255,.3) 80%,rgba(255,255,255,0) 100%)}.O0WRkf.RDPZE{-moz-box-shadow:none;box-shadow:none;color:rgba(68,68,68,0.502);cursor:default;fill:rgba(68,68,68,0.502)}.zZhnYe.RDPZE{background:rgba(153,153,153,.1)}.UxubU.RDPZE{color:rgba(255,255,255,0.502);fill:rgba(255,255,255,0.502)}.UxubU.zZhnYe.RDPZE{background:rgba(204,204,204,.1)}.CwaK9{position:relative}.RveJvd{display:inline-block;margin:.5em}.NBxL9e{-moz-transition:opacity 0.15s cubic-bezier(0.4,0,0.2,1) 0.15s;transition:opacity 0.15s cubic-bezier(0.4,0,0.2,1) 0.15s;background-color:rgba(0,0,0,.5);bottom:0;left:0;opacity:0;position:fixed;right:0;top:0;z-index:1191}.NBxL9e.iWO5td{-moz-transition:opacity 0.05s cubic-bezier(0.4,0,0.2,1);transition:opacity 0.05s cubic-bezier(0.4,0,0.2,1);opacity:1}.QSj8ac{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-orient:vertical;box-orient:vertical;flex-direction:column;bottom:0;left:0;padding:0 5%;position:absolute;right:0;top:0;transition:-webkit-transform .4s cubic-bezier(0.4,0,0.2,1);transition:transform .4s cubic-bezier(0.4,0,0.2,1);transition:transform .4s cubic-bezier(0.4,0,0.2,1),-webkit-transform .4s cubic-bezier(0.4,0,0.2,1)}.bJHJLe,.C40Us{display:block;height:3em}.pdYghb>.bJHJLe,.pdYghb>.C40Us{box-flex:1;flex-grow:1}.Inn9w{flex-shrink:1;max-height:100%}.Inn9w:focus{outline:none}.I7OXgf{-moz-box-align:stretch;box-align:stretch;align-items:stretch;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-orient:vertical;box-orient:vertical;flex-direction:column;box-shadow:0 1px 3px 0 rgba(60,64,67,.3),0 4px 8px 3px rgba(60,64,67,.15);background-color:#fff;-moz-border-radius:8px;border-radius:8px;max-width:24em;outline:1px solid transparent;overflow:hidden;position:relative;transition:-webkit-transform .225s cubic-bezier(0,0,0.2,1);transition:transform .225s cubic-bezier(0,0,0.2,1);transition:transform .225s cubic-bezier(0,0,0.2,1),-webkit-transform .225s cubic-bezier(0,0,0.2,1)}.I7OXgf.GKheFe{max-width:100%;width:400px}.I7OXgf.TcAFyb{max-width:100%;width:544px}.xiutKc .I7OXgf{padding:0}.I7OXgf.kdCdqc{transition:-webkit-transform .15s cubic-bezier(0.4,0,1,1);transition:transform .15s cubic-bezier(0.4,0,1,1);transition:transform .15s cubic-bezier(0.4,0,1,1),-webkit-transform .15s cubic-bezier(0.4,0,1,1)}.ZEeHrd.CAwICe{transform:scale(0.8)}.ZEeHrd.kdCdqc{transform:scale(0.9)}.xiutKc{-moz-box-align:stretch;box-align:stretch;align-items:stretch;padding:0}.xiutKc>.I7OXgf{box-flex:2;flex-grow:2;-moz-border-radius:0;border-radius:0;left:0;max-width:100%;right:0}.xiutKc>.C40Us,.xiutKc>.bJHJLe{box-flex:0;flex-grow:0;height:0}.df5yGe{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;flex-shrink:0;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:16px;font-weight:500;letter-spacing:.1px;line-height:24px}.VhQQpd .df5yGe{padding-bottom:0}.xiutKc .df5yGe{display:none}.feojCc{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:16px;font-weight:500;letter-spacing:.1px;line-height:24px;flex-shrink:0;box-pack:justify;justify-content:space-between;background-color:#fff;border-bottom:#dadce0 1px solid;color:#3c4043;display:none}.xiutKc .feojCc{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex}.Shk6y{box-flex:1;flex-grow:1;flex-shrink:1;margin:18px 24px 16px 24px;min-width:0;word-wrap:break-word}.Shk6y.Gx4dqb{text-align:center}.feojCc .Shk6y{margin:16px}.feojCc .Shk6y.irNx2b{margin-left:0}.feojCc .b9xlif{display:none}.jFptUc{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.df5yGe .jFptUc{display:none}.NFUcsb .ORmQmd{float:right;margin-right:4px;margin-top:4px}.UYUfn{box-flex:2;flex-grow:2;flex-shrink:2;font-family:Roboto,Arial,sans-serif;font-size:14px;font-weight:400;letter-spacing:.2px;line-height:20px;display:block;outline:none;overflow-y:auto;padding:0 24px}.fNxzgd .UYUfn{padding-top:20px}.Niudaf .UYUfn{padding-bottom:24px}.xiutKc .UYUfn{padding:16px}.OE6hId{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;flex-shrink:0;box-pack:end;justify-content:flex-end;line-height:0;padding:16px 8px 8px 24px}.xiutKc .OE6hId{display:none}.jzUkrb{box-pack:end;justify-content:flex-end;display:none}.xiutKc .jzUkrb{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;margin:0 16px}.ARrCac.O0WRkf.C0oVfc,.OE6hId .O0WRkf.C0oVfc{min-width:64px}.ARrCac+.ARrCac{margin-left:8px}.feojCc .ORmQmd{align-self:center;margin:0 4px;position:initial}.iOct6d{margin-top:8px}.hvREyb{-moz-box-align:center;align-items:center;display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-pack:center;justify-content:center}.VnX4Cd .wnIM7,.VnX4Cd .XGSlvc{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1;box-flex:1;flex-grow:1;min-width:0}.p0oLxb{transition:box-shadow 280ms cubic-bezier(0.4,0,0.2,1);-moz-user-select:none;-moz-transition:background .2s .1s;transition:background .2s .1s;border:0;-moz-border-radius:4px;border-radius:4px;color:#5f6368;cursor:pointer;display:inline-block;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:14px;font-weight:500;letter-spacing:.25px;line-height:36px;text-decoration:none;text-transform:none;min-width:auto;max-width:100%;outline:none;overflow:hidden;position:relative;text-align:center;z-index:0}.p0oLxb.iWO5td{transition:box-shadow 280ms cubic-bezier(0.4,0,0.2,1)}.p0oLxb.REtOWc{width:100%}.REtOWc .GcVcmc{justify-content:center}.CMZlRd{color:#e8eaed;fill:#e8eaed}.BEAGS{border:1px #e8eaed solid;box-sizing:border-box;color:#1a73e8;height:36px;line-height:34px}.BEAGS.iWO5td{box-shadow:0 2px 1px -1px rgba(26,115,232,0.2),0 1px 1px 0 rgba(26,115,232,0.141),0 1px 3px 0 rgba(26,115,232,0.122);border:none}.K2V86d{box-shadow:0 2px 1px -1px rgba(0,0,0,0.2),0 1px 1px 0 rgba(0,0,0,0.141),0 1px 3px 0 rgba(0,0,0,0.122);background-color:#fff;color:#1a73e8}.QkA63b{background:#1a73e8;color:#fff}.DqwBN{color:#1a73e8}.K2V86d.iWO5td{box-shadow:0 3px 5px -1px rgba(0,0,0,0.2),0 6px 10px 0 rgba(0,0,0,0.141),0 1px 18px 0 rgba(0,0,0,0.122)}.p0oLxb.QkA63b.iWO5td{box-shadow:0 3px 5px -1px rgba(26,115,232,0.2),0 6px 10px 0 rgba(26,115,232,0.141),0 1px 18px 0 rgba(26,115,232,0.122)}.GJYBjd{position:absolute;top:0;right:0;bottom:0;left:0;background-color:#5f6368;opacity:0}.CMZlRd .GJYBjd{background-color:#e8eaed}.QkA63b .GJYBjd{background-color:#fff}.DqwBN .GJYBjd,.BEAGS .GJYBjd,.K2V86d .GJYBjd{background-color:#4285f4}.p0oLxb:hover .GJYBjd{opacity:0.04}.BEAGS:hover{border-color:#d2e3fc}.QkA63b:hover{box-shadow:0 2px 1px -1px rgba(26,115,232,0.2),0 1px 1px 0 rgba(26,115,232,0.141),0 1px 3px 0 rgba(26,115,232,0.122)}.CMZlRd:hover .GJYBjd{opacity:0.04}.QkA63b:hover .GJYBjd{opacity:0.08}.p0oLxb.u3bW4e .GJYBjd{opacity:0.12}.BEAGS.u3bW4e{border-color:#d2e3fc}.CMZlRd.u3bW4e .GJYBjd{opacity:0.12}.QkA63b.u3bW4e .GJYBjd{opacity:0.24}.p0oLxb.u3bW4e:hover .GJYBjd{opacity:0.155}.CMZlRd.u3bW4e:hover .GJYBjd{opacity:0.155}.QkA63b.u3bW4e:hover .GJYBjd{opacity:0.3}.p0oLxb.RDPZE .GJYBjd{opacity:0}.bnqxkd{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,-webkit-transform 0s ease .2s;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.p0oLxb.iWO5td>.bnqxkd{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1);-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.p0oLxb.j7nIZb>.bnqxkd{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);visibility:visible}.p0oLxb>.bnqxkd{background-image:radial-gradient(circle farthest-side,rgba(0,0,0,.12),rgba(0,0,0,.12) 80%,rgba(0,0,0,0) 100%)}.CMZlRd.iWO5td>.bnqxkd{background-image:radial-gradient(circle farthest-side,rgba(255,255,255,0.161),rgba(255,255,255,0.161) 80%,rgba(255,255,255,0) 100%)}.QkA63b.iWO5td>.bnqxkd{background-image:radial-gradient(circle farthest-side,rgba(255,255,255,0.322),rgba(255,255,255,0.322) 80%,rgba(255,255,255,0) 100%)}.DqwBN.iWO5td>.bnqxkd,.BEAGS.iWO5td>.bnqxkd,.K2V86d.iWO5td>.bnqxkd{background-image:radial-gradient(circle farthest-side,rgba(66,133,244,0.161),rgba(66,133,244,0.161) 80%,rgba(66,133,244,0) 100%)}.p0oLxb.RDPZE{-moz-box-shadow:none;box-shadow:none;color:rgba(0,0,0,.38);cursor:default;fill:rgba(0,0,0,.38)}.CMZlRd.RDPZE{color:rgba(255,255,255,.38);fill:rgba(255,255,255,.38)}.BEAGS.RDPZE,.BEAGS.RDPZE:hover{border-color:rgba(0,0,0,.12)}.QkA63b.RDPZE,.K2V86d.RDPZE{background:rgba(0,0,0,.12)}.GcVcmc{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;position:relative}.GcVcmc .RdyDwe{display:inline-block;margin:0;overflow:hidden}.I0YiR .GcVcmc,.DqwBN .GcVcmc{padding:0 8px}.BEAGS .GcVcmc{padding:0 23px}.BEAGS.iWO5td .GcVcmc{padding:1px 24px}.BEAGS.iWO5td .cd29Sd.GcVcmc{padding:1px 16px 1px 12px}.BEAGS.iWO5td .rbRww.GcVcmc{padding:1px 12px 1px 16px}.BEAGS .cd29Sd.GcVcmc{padding-right:15px;padding-left:11px}.BEAGS .rbRww.GcVcmc{padding-left:15px;padding-right:11px}.QkA63b .GcVcmc,.K2V86d .GcVcmc{padding:0 24px}.GcVcmc.cd29Sd{padding:0 16px 0 12px}.GcVcmc.rbRww{padding:0 12px 0 16px}.lRRqZc{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;color:currentcolor;fill:currentcolor;margin-right:8px}.oPP9ge{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;color:currentcolor;fill:currentcolor;margin-left:8px}.JRtysb{-moz-user-select:none;-moz-transition:background .3s;transition:background .3s;border:0;-moz-border-radius:50%;border-radius:50%;color:#444;cursor:pointer;display:inline-block;fill:#444;flex-shrink:0;height:48px;outline:none;overflow:hidden;position:relative;text-align:center;width:48px;z-index:0}.JRtysb.RDPZE{cursor:default}.ZDSs1{color:rgba(255,255,255,.75);fill:rgba(255,255,255,.75)}.WzwrXb.u3bW4e{background-color:rgba(153,153,153,.4)}.ZDSs1.u3bW4e{background-color:rgba(204,204,204,.25)}.NWlf3e{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);-moz-transition:opacity .2s ease;transition:opacity .2s ease;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.JRtysb.iWO5td>.NWlf3e{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.JRtysb.j7nIZb>.NWlf3e{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);visibility:visible}.WzwrXb.iWO5td>.NWlf3e{background-image:radial-gradient(circle farthest-side,rgba(153,153,153,.4),rgba(153,153,153,.4) 80%,rgba(153,153,153,0) 100%)}.ZDSs1.iWO5td>.NWlf3e{background-image:radial-gradient(circle farthest-side,rgba(204,204,204,.25),rgba(204,204,204,.25) 80%,rgba(204,204,204,0) 100%)}.WzwrXb.RDPZE{color:rgba(68,68,68,0.502);fill:rgba(68,68,68,0.502)}.ZDSs1.RDPZE{color:rgba(255,255,255,0.502);fill:rgba(255,255,255,0.502)}.MhXXcc{line-height:44px;position:relative}.Lw7GHd{margin:8px;display:inline-block}.I12f0b:hover{background-color:rgba(32,33,36,0.039)}.I12f0b.RDPZE:hover{background-color:transparent}.hvvWV:hover{background-color:rgba(232,234,237,0.039)}.wwnMtb:hover{background-color:rgba(66,133,244,0.039)}.K2mXPb{color:#5f6368;fill:#5f6368}.hvvWV{color:#e8eaed;fill:#e8eaed}.wwnMtb{color:#1a73e8;fill:#1a73e8}.K2mXPb.u3bW4e{background-color:rgba(32,33,36,0.122)}.K2mXPb.u3bW4e:hover{background-color:rgba(32,33,36,0.157)}.hvvWV.u3bW4e{background-color:rgba(232,234,237,0.122)}.hvvWV.u3bW4e:hover{background-color:rgba(232,234,237,0.157)}.wwnMtb.u3bW4e{background-color:rgba(66,133,244,0.122)}.wwnMtb.u3bW4e:hover{background-color:rgba(66,133,244,0.157)}.I12f0b.RDPZE{color:#9aa0a6;fill:#9aa0a6}.hvvWV.RDPZE{color:rgba(255,255,255,.38);fill:rgba(255,255,255,.38)}.I12f0b .oJeWuf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:100%;width:100%}.I12f0b .snByac{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:1;flex-grow:1;justify-content:center;margin:0}.JPdR6b{-moz-transform:translateZ(0);transform:translateZ(0);-moz-transition:max-width 0.2s cubic-bezier(0,0,0.2,1),max-height 0.2s cubic-bezier(0,0,0.2,1),opacity 0.1s linear;transition:max-width 0.2s cubic-bezier(0,0,0.2,1),max-height 0.2s cubic-bezier(0,0,0.2,1),opacity 0.1s linear;background:#fff;border:0;-moz-border-radius:2px;border-radius:2px;-moz-box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);-moz-box-sizing:border-box;box-sizing:border-box;max-height:100%;max-width:100%;opacity:1;outline:1px solid transparent;z-index:2000}.XvhY1d{overflow-x:hidden;overflow-y:auto}.JAPqpe{float:left;padding:16px 0}.JPdR6b.qjTEB{-moz-transition:left 0.2s cubic-bezier(0,0,0.2,1),max-width 0.2s cubic-bezier(0,0,0.2,1),max-height 0.2s cubic-bezier(0,0,0.2,1),opacity 0.05s linear,top 0.2s cubic-bezier(0,0,0.2,1);transition:left 0.2s cubic-bezier(0,0,0.2,1),max-width 0.2s cubic-bezier(0,0,0.2,1),max-height 0.2s cubic-bezier(0,0,0.2,1),opacity 0.05s linear,top 0.2s cubic-bezier(0,0,0.2,1)}.JPdR6b.jVwmLb{max-height:56px;opacity:0}.JPdR6b.CAwICe{overflow:hidden}.JPdR6b.oXxKqf{-moz-transition:none;transition:none}.z80M1{color:#222;cursor:pointer;display:block;outline:none;overflow:hidden;padding:0 24px;position:relative}.uyYuVb{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;font-size:14px;font-weight:400;line-height:40px;height:40px;position:relative;white-space:nowrap}.jO7h3c{box-flex:1;flex-grow:1;min-width:0}.JPdR6b.e5Emjc .z80M1{padding-left:64px}.JPdR6b.CblTmf .z80M1{padding-right:48px}.PCdOIb{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;flex-direction:column;justify-content:center;background-repeat:no-repeat;height:40px;left:24px;opacity:0.54;position:absolute}.z80M1.RDPZE .PCdOIb{opacity:0.26}.z80M1.FwR7Pc{outline:1px solid transparent;background-color:#eee}.z80M1.RDPZE{color:#b8b8b8;cursor:default}.z80M1.N2RpBe::before{-moz-transform:rotate(45deg);transform:rotate(45deg);-moz-transform-origin:left;transform-origin:left;content:"\0000a0";display:block;border-right:2px solid #222;border-bottom:2px solid #222;height:16px;left:24px;opacity:0.54;position:absolute;top:13%;width:7px;z-index:0}.JPdR6b.CblTmf .z80M1.N2RpBe::before{left:auto;right:16px}.z80M1.RDPZE::before{border-color:#b8b8b8;opacity:1}.aBBjbd{pointer-events:none;position:absolute}.z80M1.qs41qe>.aBBjbd{-moz-animation:quantumWizBoxInkSpread 0.3s ease-out;animation:quantumWizBoxInkSpread 0.3s ease-out;animation-fill-mode:forwards;background-image:-moz-radial-gradient(circle farthest-side,#bdbdbd,#bdbdbd 80%,rgba(189,189,189,0) 100%);background-image:radial-gradient(circle farthest-side,#bdbdbd,#bdbdbd 80%,rgba(189,189,189,0) 100%);background-size:cover;opacity:1;top:0;left:0}.J0XlZe{color:inherit;line-height:40px;padding:0 6px 0 1em}.a9caSc{color:inherit;direction:ltr;padding:0 6px 0 1em}.kCtYwe{border-top:1px solid rgba(0,0,0,.12);margin:7px 0}.B2l7lc{border-left:1px solid rgba(0,0,0,.12);display:inline-block;height:48px}@media screen and (max-width:840px){.JAPqpe{padding:8px 0}.z80M1{padding:0 16px}.JPdR6b.e5Emjc .z80M1{padding-left:48px}.PCdOIb{left:12px}}.jgvuAb{-moz-user-select:none;-moz-transition:background .3s;transition:background .3s;border:0;-moz-border-radius:3px;border-radius:3px;color:#444;cursor:pointer;display:inline-block;font-size:14px;font-weight:500;outline:none;position:relative;text-align:center}.jgvuAb.u3bW4e{background-color:rgba(153,153,153,.4)}.kRoyt{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);transition:-webkit-transform 0 linear .2s,opacity .2s ease;transition:opacity .2s ease,-webkit-transform 0 linear .2s;transition:transform 0 linear .2s,opacity .2s ease;transition:transform 0 linear .2s,opacity .2s ease,-webkit-transform 0 linear .2s;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.jgvuAb.qs41qe .ziS7vd{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.jgvuAb .kRoyt{background-image:radial-gradient(circle farthest-side,rgba(153,153,153,.4),rgba(153,153,153,.4) 80%,rgba(153,153,153,0) 100%)}.jgvuAb.RDPZE{-moz-box-shadow:none;box-shadow:none;color:rgba(68,68,68,0.502);cursor:default}.vRMGwf{position:relative}.e2CuFe{border-color:rgba(68,68,68,.4) transparent;border-style:solid;border-width:6px 6px 0 6px;height:0;width:0;position:absolute;right:5px;top:15px}.CeEBt{position:absolute;right:0;top:0;width:24px;overflow:hidden}.ncFHed{-moz-transition:opacity 0.1s linear;transition:opacity 0.1s linear;background:#fff;border:0;-moz-box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);opacity:0;outline:1px solid transparent;overflow:hidden;overflow-y:auto;position:fixed;z-index:2000}.jgvuAb.iWO5td .ncFHed{opacity:1}.MocG8c{border-color:transparent;color:#222;height:0;list-style:none;outline:none;overflow:hidden;padding-left:16px;padding-right:24px;position:relative;text-align:left;white-space:nowrap}.MocG8c.RDPZE{color:#b8b8b8;pointer-events:none;cursor:default}.MocG8c.DEh1R{color:rgba(0,0,0,.54)}.jgvuAb.e5Emjc .MocG8c{padding-left:48px}.ry3kXd .MocG8c.KKjvXb{height:auto;padding-bottom:8px;padding-top:8px}.Ulgu9 .MocG8c:not(.KKjvXb){width:0;border:0;margin:0;position:relative;opacity:.0001;padding:0;top:-99999px;pointer-events:none}.ncFHed .MocG8c{cursor:pointer;height:auto;padding-right:26px;padding-bottom:8px;padding-top:8px}.ncFHed .MocG8c.KKjvXb{background-color:#eee;border-style:dotted;border-width:1px 0;outline:1px solid transparent;padding-bottom:7px;padding-top:7px}.MWQFLe{background-repeat:no-repeat;height:21px;left:12px;opacity:0.54;position:absolute;right:auto;top:5px;vertical-align:middle;width:21px}.ncFHed .MocG8c.KKjvXb .MWQFLe{top:4px}.jgvuAb.RDPZE .MWQFLe,.MocG8c.RDPZE .MWQFLe{opacity:0.26}.ncFHed.qs41qe .ziS7vd{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.VOUU9e{border-top:0;height:0;margin:0;overflow:hidden}.ncFHed .VOUU9e{border-top:1px solid rgba(0,0,0,.12);margin:7px 0}.mAW2Ib{width:64px}.YuHtjc .KKjvXb .vRMGwf{visibility:hidden}.YuHtjc .MocG8c{padding-left:48px;padding-right:12px}.ybOdnf .oJeWuf{line-height:32px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;overflow:hidden}.ybOdnf .eU809d{top:22px;right:19px;border-color:#5f6368 transparent;border-width:5px 5px 0 5px}.ybOdnf.iWO5td .eU809d{transform:scaleY(-1);border-color:#bdc1c6 transparent}.ybOdnf:not(.iWO5td) .LMgvRb.KKjvXb{-moz-border-radius:4px;border-radius:4px}.ybOdnf .OA0qNb{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);padding:8px 0 8px 0;-moz-border-radius:4px;border-radius:4px}.cr8auc{background-color:#f8f9fa}.ybOdnf.iWO5td{background-color:#e8f0fe}.ybOdnf .OA0qNb .LMgvRb[aria-selected="true"]{background-color:rgba(26,115,232,0.078)}.ybOdnf .OA0qNb .LMgvRb[aria-selected="true"]:hover{background-color:rgba(26,115,232,0.039)}.HZ3kWc{font-family:Roboto,Arial,sans-serif;font-size:14px;font-weight:400;letter-spacing:.2px;line-height:20px;color:#202124;max-width:280px;min-width:112px;padding-right:48px}.RDPZE .HZ3kWc{color:rgba(0,0,0,.38)}.ybOdnf.llrsB .HZ3kWc{max-width:none}.HZ3kWc .uLX2p{height:24px;opacity:1;top:12px;width:24px}.HZ3kWc.KKjvXb .uLX2p.uLX2p{top:11px}.mbHMhf{border-top:0;height:0;margin:0;overflow:hidden}.QXL7Te .mbHMhf{border-top:1px solid rgba(0,0,0,.12);margin:8px 0}@keyframes agmTextInputRemoveUnderline{0%{-moz-transform:scaleX(1);transform:scaleX(1);opacity:1}to{-moz-transform:scaleX(1);transform:scaleX(1);opacity:0}}@keyframes agmTextInputAddUnderline{0%{-moz-transform:scaleX(0);transform:scaleX(0)}to{-moz-transform:scaleX(1);transform:scaleX(1)}}.W9wDc{-moz-user-select:none;-moz-user-select:none;display:inline-block;outline:none;width:280px}.W9wDc.YcPWMc{width:100%}.n9IS1{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-align:center;box-align:center;align-items:center;position:relative}.W9wDc.F5VHze .n9IS1,.W9wDc.F5VHze .FtBNWb{-moz-box-orient:horizontal;-moz-box-direction:reverse;flex-direction:row-reverse}.HyS0Qd .n9IS1{background-color:#f8f9fa;-moz-border-radius:4px 4px 0 0;border-radius:4px 4px 0 0;height:56px}.HyS0Qd.RDPZE .n9IS1{background-color:rgba(248,249,250,.38)}.HyS0Qd:not(.RDPZE):hover .n9IS1{background-color:#f1f3f4;cursor:pointer}.D3oBEe .n9IS1:before{-moz-border-radius:4px;border-radius:4px;border:1px solid #dadce0;bottom:0;content:"";left:0;position:absolute;right:0;top:0;z-index:0}.D3oBEe.u3bW4e .n9IS1:before{border:2px solid #1a73e8}.D3oBEe.IYewr .n9IS1:before{border:2px solid #d93025}.D3oBEe.IYewr.RDPZE .n9IS1:before{border-color:rgba(217,48,37,.38)}.FtBNWb{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;box-flex:1;flex-grow:1;flex-shrink:1;cursor:text;min-width:0%;position:relative}.poFWNe{box-flex:1;flex-grow:1;flex-shrink:1;font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;background-color:transparent;border:none;-moz-box-sizing:content-box;box-sizing:content-box;caret-color:#1a73e8;display:block;height:24px;margin:0;padding:16px;min-width:0%;outline:none;z-index:0}.poFWNe[disabled]{color:rgba(60,64,67,.38)}.HyS0Qd:not(.yaevDc) .poFWNe{padding:23px 16px 9px 16px}.poFWNe:invalid,.poFWNe:-moz-submit-invalid,.poFWNe:-moz-ui-invalid{-moz-box-shadow:none;box-shadow:none}.W9wDc.HYyP9e .poFWNe{padding-left:0}.W9wDc.JFSSzd .poFWNe{padding-left:4px}.W9wDc.svmwUe:not(.F5VHze) .poFWNe{padding-right:0}.W9wDc.svmwUe.F5VHze .poFWNe{padding-right:0}.W9wDc.vkREqc:not(.F5VHze) .poFWNe{padding-right:4px}.W9wDc.vkREqc.F5VHze .poFWNe{padding-right:4px}.W9wDc.IYewr .poFWNe{caret-color:#d93025}.rXTzdc .poFWNe::-ms-clear,.rXTzdc .poFWNe::-ms-reveal{display:none}.CROdRc+.poFWNe{padding-left:2px}.AKIybd{background-color:#80868b;bottom:0;height:1px;left:0;margin:0;padding:0;position:absolute;width:100%}.AKIybd:before{content:"";position:absolute;top:0;bottom:-1px;left:0;right:0;border-bottom:1px solid rgba(0,0,0,0);pointer-events:none}.HyS0Qd.RDPZE .AKIybd{background-color:rgba(128,134,139,.38)}.cWL65e{-moz-transform:scaleX(0);transform:scaleX(0);background-color:#1a73e8;bottom:0;height:2px;left:0;margin:0;padding:0;position:absolute;width:100%}.D3oBEe .AKIybd,.D3oBEe .cWL65e{display:none}.W9wDc.IYewr .AKIybd,.W9wDc.IYewr .cWL65e{background-color:#d93025;height:2px}.W9wDc.IYewr.RDPZE .AKIybd,.W9wDc.IYewr.RDPZE .cWL65e{background-color:rgba(217,48,37,.38)}.poFWNe[disabled]~.AKIybd{background:none;border-bottom:1px dotted #dadce0}.cWL65e.Y2Zypf{-moz-animation:agmTextInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:agmTextInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1)}.W9wDc.u3bW4e .cWL65e{-moz-animation:agmTextInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:agmTextInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);-moz-transform:scaleX(1);transform:scaleX(1)}.qTs5Xc{-moz-transform-origin:bottom left;transform-origin:bottom left;-moz-transition:all .3s cubic-bezier(0.4,0,0.2,1);transition:all .3s cubic-bezier(0.4,0,0.2,1);transition-property:color,-webkit-transform;transition-property:color,transform;transition-property:color,transform,-webkit-transform;font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;color:#5f6368;left:16px;right:16px;text-overflow:ellipsis;overflow:hidden;white-space:nowrap;pointer-events:none;position:absolute;top:16px}.D3oBEe .qTs5Xc{background-color:white;left:12px;max-width:-moz-calc(100% - 32px);max-width:calc(100% - 32px);padding:2px 4px;right:auto;top:14px}.D3oBEe .poFWNe:not([disabled]):focus~.qTs5Xc,.D3oBEe .poFWNe[badinput=true]~.qTs5Xc,.W9wDc.D3oBEe.CDELXb .qTs5Xc,.W9wDc.D3oBEe.sM9l1e .qTs5Xc{-moz-transform:scale(.75) translateY(-41px);transform:scale(.75) translateY(-41px)}.W9wDc.RDPZE .qTs5Xc{color:rgba(60,64,67,.38)}.W9wDc.HYyP9e .qTs5Xc{left:0}.D3oBEe .n9IS1>.qTs5Xc{left:12px}.HyS0Qd.svmwUe .qTs5Xc{right:0}.poFWNe:not([disabled]):focus~.qTs5Xc,.poFWNe[badinput=true]~.qTs5Xc,.W9wDc.CDELXb .qTs5Xc,.W9wDc.sM9l1e .qTs5Xc{-moz-transform:scale(.75) translateY(-20px);transform:scale(.75) translateY(-20px)}.poFWNe:not([disabled]):focus~.qTs5Xc{color:#1a73e8}.W9wDc.IYewr .poFWNe:not([disabled]):focus~.qTs5Xc,.W9wDc.IYewr .n9IS1 .qTs5Xc{color:#d93025}.W9wDc.IYewr.RDPZE .n9IS1 .qTs5Xc{color:rgba(217,48,37,.38)}.uUUR3b{font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;color:#9aa0a6;left:16px;overflow:hidden;pointer-events:none;position:absolute;right:16px;text-overflow:ellipsis;top:16px;white-space:nowrap}.W9wDc.RDPZE .uUUR3b{color:rgba(154,160,166,.38)}.HyS0Qd:not(.yaevDc) .uUUR3b{top:23px}.W9wDc.CDELXb .uUUR3b{display:none}.W9wDc.HYyP9e .uUUR3b{left:0}.W9wDc.svmwUe .uUUR3b{right:0}.uDjDl{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex}.DAKCob{font-family:Roboto,Arial,sans-serif;font-size:12px;font-weight:400;letter-spacing:.3px;line-height:16px;height:16px;margin-left:auto;padding:4px 12px;pointer-events:none;white-space:nowrap}.uNeeU,.cHUCT:not(:empty){flex:1 1 auto;font-family:Roboto,Arial,sans-serif;font-size:12px;font-weight:400;letter-spacing:.3px;line-height:16px;min-height:16px;padding:4px 16px}.cHUCT{pointer-events:none}.uNeeU{color:#d93025}.W9wDc.RDPZE .uNeeU{color:rgba(217,48,37,.38)}.cHUCT,.DAKCob{color:#5f6368}.W9wDc.RDPZE .cHUCT,.W9wDc.RDPZE .DAKCob{color:rgba(95,99,104,.38)}.W9wDc.IYewr .cHUCT,.W9wDc:not(.IYewr) .cHUCT:not(:empty)+.uNeeU{display:none}.hmzrif,.Hzgwd{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;box-flex:0;flex-grow:0;flex-shrink:0;font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;align-self:center;color:#80868b;height:24px}.W9wDc.svmwUe:not(.F5VHze) .n9IS1 .hmzrif{padding-right:0}.W9wDc.svmwUe.F5VHze .n9IS1 .hmzrif{padding-right:0}.W9wDc.HYyP9e:not(.F5VHze) .n9IS1 .Hzgwd{padding-left:0}.W9wDc.HYyP9e.F5VHze .n9IS1 .Hzgwd{padding-left:0}.W9wDc.RDPZE .hmzrif,.W9wDc.RDPZE .Hzgwd{opacity:.38}.W9wDc:not(.F5VHze) .hmzrif{padding:16px 16px 16px 0}.W9wDc.F5VHze .hmzrif{padding:16px 16px 16px 0}.W9wDc:not(.F5VHze) .Hzgwd{padding:16px 0 16px 16px}.W9wDc.F5VHze .Hzgwd{padding:16px 0 16px 16px}.HyS0Qd:not(.yaevDc):not(.F5VHze) .hmzrif{padding:24px 16px 8px 0}.HyS0Qd:not(.yaevDc).F5VHze .hmzrif{padding:24px 16px 8px 0}.HyS0Qd:not(.yaevDc):not(.F5VHze) .Hzgwd{padding:24px 0 8px 16px}.HyS0Qd:not(.yaevDc).F5VHze .Hzgwd{padding:24px 0 8px 16px}.Pl5mpf,.GIwIzd{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-sizing:border-box;box-sizing:border-box;height:100%;line-height:24px;padding:0 12px;position:relative}.CROdRc{align-self:center;padding:16px 0 16px 16px}.HyS0Qd:not(.yaevDc) .CROdRc{padding:23px 0 9px 16px}.ndfHFb-c4YZDc-K9a4Re{position:absolute;-moz-transition:bottom .218s ease-out;transition:bottom .218s ease-out;left:0;right:0;top:0;bottom:0;z-index:0}.fFW7wc-L5Fo6c.fFW7wc-jJNx8e{-moz-box-shadow:rgba(0,0,0,.2) 0 4px 16px;-moz-box-shadow:rgba(0,0,0,.2) 0 4px 16px;box-shadow:rgba(0,0,0,.2) 0 4px 16px;color:#000;padding:0;position:absolute;z-index:1002}.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-OEVmcd-yHKmmc{background-color:#f1f1f1}.fFW7wc-L5Fo6c.fFW7wc-HLvlvd-Hn6s1b.fFW7wc-VWkKje .fFW7wc-jJNx8e-OEVmcd-yHKmmc{background-color:#fff}.fFW7wc-L5Fo6c.fFW7wc-jJNx8e.VIpgJd-xl07Ob{border-color:#ccc;line-height:0;max-height:none;overflow:visible}.fFW7wc-L5Fo6c.fFW7wc-jJNx8e-ma6Yeb{margin-top:15px}.fFW7wc-L5Fo6c.fFW7wc-VWkKje.fFW7wc-jJNx8e-ma6Yeb{margin-top:9px}.fFW7wc-L5Fo6c.fFW7wc-jJNx8e-cGMI2b{margin-top:-15px}.fFW7wc-L5Fo6c.fFW7wc-VWkKje.fFW7wc-jJNx8e-cGMI2b{margin-top:-9px}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc,.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW{position:absolute;width:32px;z-index:0}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc{top:-15px}.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-yHKmmc{top:-10px;width:20px}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW{bottom:-16px}.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-hgHJW{bottom:-10px;width:20px}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-SmKAyb,.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-VtOx3e{border:16px solid;height:0;position:absolute;width:0}.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-SmKAyb,.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-VtOx3e{border:10px solid}.fFW7wc-L5Fo6c.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb{border-color:#f1f1f1 transparent}.fFW7wc-L5Fo6c.fFW7wc-HLvlvd-Hn6s1b.fFW7wc-VWkKje .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb{border-color:#fff transparent}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb{border-color:#fff transparent;top:1px;z-index:1}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-SmKAyb{border-color:#fff transparent;bottom:1px;z-index:1}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-VtOx3e{border-color:rgba(0,0,0,.2) transparent}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-VtOx3e{border-color:rgba(0,0,0,.2) transparent;bottom:0}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-SmKAyb,.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-yHKmmc .fFW7wc-jJNx8e-hFsbo-VtOx3e{border-top-width:0}.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-SmKAyb,.fFW7wc-L5Fo6c .fFW7wc-jJNx8e-hFsbo-hgHJW .fFW7wc-jJNx8e-hFsbo-VtOx3e{border-bottom-width:0}.ndfHFb-c4YZDc{color:#fff;font-family:arial,sans-serif;overflow:clip;opacity:0;visibility:hidden;-moz-transition-property:opacity,visibility;transition-property:opacity,visibility;-moz-transition-duration:0.1s,0s;transition-duration:0.1s,0s;-moz-transition-timing-function:cubic-bezier(0,0,0.2,1);transition-timing-function:cubic-bezier(0,0,0.2,1);-moz-transition-delay:0s,0.1s;transition-delay:0s,0.1s;position:fixed;top:0;bottom:0;left:0;right:0;z-index:1193}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb{font-family:"Google Sans",Roboto,arial,sans-serif}.ndfHFb-c4YZDc-TSZdd{opacity:1;visibility:visible;-moz-transition-timing-function:cubic-bezier(0.4,0,1,1);transition-timing-function:cubic-bezier(0.4,0,1,1);-moz-transition-delay:0s,0s;transition-delay:0s,0s}.ndfHFb-c4YZDc-bnBfGc{background-color:#1e1e1e;position:fixed;top:0;bottom:0;left:0;right:0;filter:alpha(opacity=93);opacity:.93}.ndfHFb-c4YZDc-JNEHMb{left:0;position:absolute;right:0}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-bnBfGc{background-color:#d1d1d1;filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-bnBfGc{background-color:rgba(0,0,0,.85);filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-bnBfGc{background-color:rgba(31,31,31,.92)}.ndfHFb-c4YZDc-qbOKL-OEVmcd{margin:0;height:100%;width:100%;overflow:hidden!important}.ndfHFb-c4YZDc-AHmuwe-Hr88gd-OWB6Me *:focus{outline:none}.VIpgJd-TzA9Ye-eEGnhe{position:relative;display:-moz-inline-box;display:inline-block}* html .VIpgJd-TzA9Ye-eEGnhe{display:inline}*:first-child+html .VIpgJd-TzA9Ye-eEGnhe{display:inline}.C0oVfc{line-height:20px;min-width:88px}.C0oVfc .RveJvd{margin:8px}.llhEMd{-moz-transition:opacity .15s cubic-bezier(0.4,0,0.2,1) .15s;transition:opacity .15s cubic-bezier(0.4,0,0.2,1) .15s;background-color:rgba(0,0,0,0.502);bottom:0;left:0;opacity:0;position:fixed;right:0;top:0;z-index:1191}.llhEMd.iWO5td{-moz-transition:opacity .05s cubic-bezier(0.4,0,0.2,1);transition:opacity .05s cubic-bezier(0.4,0,0.2,1);opacity:1}.mjANdc{transition:-webkit-transform .4s cubic-bezier(0.4,0,0.2,1);transition:transform .4s cubic-bezier(0.4,0,0.2,1);transition:transform .4s cubic-bezier(0.4,0,0.2,1),-webkit-transform .4s cubic-bezier(0.4,0,0.2,1);-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-orient:vertical;box-orient:vertical;flex-direction:column;bottom:0;left:0;padding:0 5%;position:absolute;right:0;top:0}.x3wWge,.ONJhl{display:block;height:3em}.eEPege>.x3wWge,.eEPege>.ONJhl{box-flex:1;flex-grow:1}.J9Nfi{flex-shrink:1;max-height:100%}.g3VIld{-moz-box-align:stretch;box-align:stretch;align-items:stretch;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-orient:vertical;box-orient:vertical;flex-direction:column;transition:-webkit-transform .225s cubic-bezier(0,0,0.2,1);transition:transform .225s cubic-bezier(0,0,0.2,1);transition:transform .225s cubic-bezier(0,0,0.2,1),-webkit-transform .225s cubic-bezier(0,0,0.2,1);position:relative;background-color:#fff;-moz-border-radius:2px;border-radius:2px;-moz-box-shadow:0 12px 15px 0 rgba(0,0,0,.24);box-shadow:0 12px 15px 0 rgba(0,0,0,.24);max-width:24em;outline:1px solid transparent;overflow:hidden}.vcug3d .g3VIld{padding:0}.g3VIld.kdCdqc{transition:-webkit-transform .15s cubic-bezier(0.4,0,1,1);transition:transform .15s cubic-bezier(0.4,0,1,1);transition:transform .15s cubic-bezier(0.4,0,1,1),-webkit-transform .15s cubic-bezier(0.4,0,1,1)}.Up8vH.CAwICe{transform:scale(0.8)}.Up8vH.kdCdqc{transform:scale(0.9)}.vcug3d{-moz-box-align:stretch;box-align:stretch;align-items:stretch;padding:0}.vcug3d>.g3VIld{box-flex:2;flex-grow:2;-moz-border-radius:0;border-radius:0;left:0;right:0;max-width:100%}.vcug3d>.ONJhl,.vcug3d>.x3wWge{box-flex:0;flex-grow:0;height:0}.tOrNgd{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;flex-shrink:0;font:500 20px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;padding:24px 24px 20px 24px}.vcug3d .tOrNgd{display:none}.TNczib{box-pack:justify;justify-content:space-between;flex-shrink:0;-moz-box-shadow:0 3px 4px 0 rgba(0,0,0,.24);box-shadow:0 3px 4px 0 rgba(0,0,0,.24);background-color:#455a64;color:white;display:none;font:500 20px Roboto,RobotoDraft,Helvetica,Arial,sans-serif}.vcug3d .TNczib{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex}.PNenzf{box-flex:1;flex-grow:1;flex-shrink:1;overflow:hidden;word-wrap:break-word}.TNczib .PNenzf{margin:16px 0}.VY7JQd{height:0}.TNczib .VY7JQd,.tOrNgd .bZWIgd{display:none}.R6Lfte .Wtw8H{flex-shrink:0;display:block;margin:-12px -6px 0 0}.PbnGhe{box-flex:2;flex-grow:2;flex-shrink:2;display:block;font:400 14px/20px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;padding:0 24px;overflow-y:auto}.Whe8ub .PbnGhe{padding-top:24px}.hFEqNb .PbnGhe{padding-bottom:24px}.vcug3d .PbnGhe{padding:16px}.XfpsVe{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;flex-shrink:0;box-pack:end;justify-content:flex-end;padding:24px 24px 16px 24px}.vcug3d .XfpsVe{display:none}.OllbWe{box-pack:end;justify-content:flex-end;display:none}.vcug3d .OllbWe{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-align:start;box-align:start;align-items:flex-start;margin:0 16px}.kHssdc.O0WRkf.C0oVfc,.XfpsVe .O0WRkf.C0oVfc{min-width:64px}.kHssdc+.kHssdc{margin-left:8px}.TNczib .kHssdc{color:#fff;margin-top:10px}.TNczib .Wtw8H{margin:4px 24px 4px 0}.TNczib .kHssdc.u3bW4e,.TNczib .Wtw8H.u3bW4e{background-color:rgba(204,204,204,.25)}.TNczib .kHssdc>.Vwe4Vb,.TNczib .Wtw8H>.VTBa7b{background-image:radial-gradient(circle farthest-side,rgba(255,255,255,.3),rgba(255,255,255,.3) 80%,rgba(255,255,255,0) 100%)}.TNczib .kHssdc.RDPZE,.TNczib .Wtw8H.RDPZE{color:rgba(255,255,255,.5);fill:rgba(255,255,255,.5)}.c7fp5b{-moz-user-select:none;-moz-transition:background .3s;transition:background .3s;border:0;-moz-border-radius:3px;border-radius:3px;color:#444;cursor:pointer;display:inline-block;font-size:14px;font-weight:500;min-width:88px;outline:none;overflow:hidden;position:relative;text-align:center}.hhcOmc{color:#fff;fill:#fff}.JvtX2e{-moz-transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);background:#dfdfdf;-moz-box-shadow:0px 2px 2px 0px rgba(0,0,0,.14),0px 3px 1px -2px rgba(0,0,0,.12),0px 1px 5px 0px rgba(0,0,0,.2);box-shadow:0px 2px 2px 0px rgba(0,0,0,.14),0px 3px 1px -2px rgba(0,0,0,.12),0px 1px 5px 0px rgba(0,0,0,.2)}.rGMe1e{background:#4285f4;color:#fff}.JvtX2e.qs41qe{-moz-transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);transition:box-shadow .28s cubic-bezier(0.4,0,0.2,1);-moz-transition:background .8s;transition:background .8s;-moz-box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2)}.rGMe1e.qs41qe{background:#3367d6}.JvtX2e.RDPZE{background:rgba(153,153,153,.1)}.g4jUVc{-moz-transition:opacity .2s ease;transition:opacity .2s ease;background-color:rgba(0,0,0,0.122);bottom:0;left:0;opacity:0;pointer-events:none;position:absolute;right:0;top:0}.FS4hgd.u3bW4e{background-color:rgba(153,153,153,.4)}.hhcOmc.u3bW4e{background-color:rgba(204,204,204,.25)}.JvtX2e.u3bW4e .g4jUVc{opacity:1}.lVYxmb{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);-moz-transition:opacity .2s ease;transition:opacity .2s ease;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0;visibility:hidden}.c7fp5b.iWO5td>.lVYxmb{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1;visibility:visible}.c7fp5b.j7nIZb>.lVYxmb{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);visibility:visible}.c7fp5b>.lVYxmb{background-image:radial-gradient(circle farthest-side,rgba(153,153,153,.4),rgba(153,153,153,.4) 80%,rgba(153,153,153,0) 100%)}.FS4hgd.iWO5td>.lVYxmb{background-image:radial-gradient(circle farthest-side,rgba(153,153,153,.4),rgba(153,153,153,.4) 80%,rgba(153,153,153,0) 100%)}.hhcOmc.iWO5td>.lVYxmb{background-image:radial-gradient(circle farthest-side,rgba(204,204,204,.25),rgba(204,204,204,.25) 80%,rgba(204,204,204,0) 100%)}.FS4hgd.RDPZE{color:rgba(68,68,68,0.502);fill:rgba(68,68,68,0.502);cursor:default}.hhcOmc.RDPZE{color:rgba(255,255,255,0.502);fill:rgba(255,255,255,0.502)}.c7fp5b.RDPZE{-moz-box-shadow:none;box-shadow:none;color:rgba(68,68,68,0.502);cursor:default}.I3EnF{position:relative;margin:16px}.NlWrkb{display:inline-block;line-height:48px}.rFrNMe{-moz-user-select:none;-moz-user-select:none;display:inline-block;outline:none;padding-bottom:8px;width:200px}.aCsJod{height:40px;position:relative;vertical-align:top}.aXBtI{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;position:relative;top:14px}.Xb9hP{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1;box-flex:1;flex-grow:1;flex-shrink:1;min-width:0%;position:relative}.A37UZe{-moz-box-sizing:border-box;box-sizing:border-box;height:24px;line-height:24px;position:relative}.qgcB3c:not(:empty){padding-right:12px}.sxyYjd:not(:empty){padding-left:12px}.whsOnd{-moz-box-flex:1;box-flex:1;flex-grow:1;flex-shrink:1;background-color:transparent;border:none;display:block;font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:24px;line-height:24px;margin:0;min-width:0%;outline:none;padding:0;z-index:0}.rFrNMe.dm7YTc .whsOnd{color:#fff}.whsOnd:invalid,.whsOnd:-moz-submit-invalid,.whsOnd:-moz-ui-invalid{-moz-box-shadow:none;box-shadow:none}.I0VJ4d>.whsOnd::-ms-clear,.I0VJ4d>.whsOnd::-ms-reveal{display:none}.i9lrp{background-color:rgba(0,0,0,.12);bottom:-2px;height:1px;left:0;margin:0;padding:0;position:absolute;width:100%}.i9lrp:before{content:"";position:absolute;top:0;bottom:-2px;left:0;right:0;border-bottom:1px solid rgba(0,0,0,0);pointer-events:none}.rFrNMe.dm7YTc .i9lrp{background-color:rgba(255,255,255,.7)}.OabDMe{transform:scaleX(0);background-color:#4285f4;bottom:-2px;height:2px;left:0;margin:0;padding:0;position:absolute;width:100%}.rFrNMe.dm7YTc .OabDMe{background-color:#a1c2fa}.rFrNMe.k0tWj .i9lrp,.rFrNMe.k0tWj .OabDMe{background-color:#d50000;height:2px}.rFrNMe.k0tWj.dm7YTc .i9lrp,.rFrNMe.k0tWj.dm7YTc .OabDMe{background-color:#e06055}.whsOnd[disabled]{color:rgba(0,0,0,.38)}.rFrNMe.dm7YTc .whsOnd[disabled]{color:rgba(255,255,255,.5)}.whsOnd[disabled]~.i9lrp{background:none;border-bottom:1px dotted rgba(0,0,0,.38)}.OabDMe.Y2Zypf{animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1)}.rFrNMe.u3bW4e .OabDMe{animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);transform:scaleX(1)}.rFrNMe.sdJrJc>.aCsJod{padding-top:24px}.AxOyFc{transform-origin:bottom left;transition:all .3s cubic-bezier(0.4,0,0.2,1);transition-property:color,bottom,-webkit-transform;transition-property:color,bottom,transform;transition-property:color,bottom,transform,-webkit-transform;color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-size:16px;pointer-events:none;position:absolute;bottom:3px;left:0;width:100%}.whsOnd:not([disabled]):focus~.AxOyFc,.whsOnd[badinput=true]~.AxOyFc,.rFrNMe.CDELXb .AxOyFc,.rFrNMe.dLgj8b .AxOyFc{transform:scale(0.75) translateY(-39px)}.whsOnd:not([disabled]):focus~.AxOyFc{color:#3367d6}.rFrNMe.dm7YTc .whsOnd:not([disabled]):focus~.AxOyFc{color:#a1c2fa}.rFrNMe.k0tWj .whsOnd:not([disabled]):focus~.AxOyFc{color:#d50000}.ndJi5d{color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;max-width:100%;overflow:hidden;pointer-events:none;position:absolute;text-overflow:ellipsis;top:2px;left:0;white-space:nowrap}.rFrNMe.CDELXb .ndJi5d{display:none}.K0Y8Se{font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:16px;margin-left:auto;padding-left:16px;padding-top:8px;pointer-events:none;opacity:.3;white-space:nowrap}.rFrNMe.dm7YTc .AxOyFc,.rFrNMe.dm7YTc .K0Y8Se,.rFrNMe.dm7YTc .ndJi5d{color:rgba(255,255,255,.7)}.rFrNMe.Tyc9J{padding-bottom:4px}.dEOOab,.ovnfwe:not(:empty){-moz-box-flex:1;-moz-box-flex:1 1 auto;flex:1 1 auto;font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;min-height:16px;padding-top:8px}.LXRPh{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.ovnfwe{pointer-events:none}.dEOOab{color:#d50000}.rFrNMe.dm7YTc .dEOOab,.rFrNMe.dm7YTc.k0tWj .whsOnd:not([disabled]):focus~.AxOyFc{color:#e06055}.ovnfwe{opacity:.3}.rFrNMe.dm7YTc .ovnfwe{color:rgba(255,255,255,.7);opacity:1}.rFrNMe.k0tWj .ovnfwe,.rFrNMe:not(.k0tWj) .ovnfwe:not(:empty)+.dEOOab{display:none}@keyframes quantumWizPaperInputRemoveUnderline{0%{transform:scaleX(1);opacity:1}to{transform:scaleX(1);opacity:0}}@keyframes quantumWizPaperInputAddUnderline{0%{transform:scaleX(0)}to{transform:scaleX(1)}}.edhGSc{-moz-user-select:none;-moz-user-select:none;display:inline-block;outline:none;padding-bottom:8px}.RpC4Ne{min-height:1.5em;position:relative;vertical-align:top}.Pc9Gce{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;position:relative;padding-top:14px}.KHxj8b{-moz-box-flex:1;box-flex:1;flex-grow:1;flex-shrink:1;background-color:transparent;border:none;display:block;font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:24px;min-height:24px;line-height:24px;margin:0;outline:none;padding:0;resize:none;white-space:pre-wrap;word-wrap:break-word;z-index:0;overflow-y:visible;overflow-x:hidden}.KHxj8b.VhWN2c{text-align:center}.edhGSc.dm7YTc .KHxj8b{color:rgba(255,255,255,.87)}.edhGSc.u3bW4e.dm7YTc .KHxj8b{color:#fff}.z0oSpf{background-color:rgba(0,0,0,.12);height:1px;left:0;margin:0;padding:0;position:absolute;width:100%}.edhGSc.dm7YTc>.RpC4Ne>.z0oSpf{background-color:rgba(255,255,255,.12)}.Bfurwb{transform:scaleX(0);background-color:#4285f4;height:2px;left:0;margin:0;padding:0;position:absolute;width:100%}.edhGSc.k0tWj>.RpC4Ne>.z0oSpf,.edhGSc.k0tWj>.RpC4Ne>.Bfurwb{background-color:#d50000;height:2px}.edhGSc.k0tWj.dm7YTc>.RpC4Ne>.z0oSpf,.edhGSc.k0tWj.dm7YTc>.RpC4Ne>.Bfurwb{background-color:#ff6e6e}.edhGSc.RDPZE .KHxj8b{color:rgba(0,0,0,.38)}.edhGSc.RDPZE>.RpC4Ne>.z0oSpf{background:none;border-bottom:1px dotted rgba(0,0,0,.38)}.Bfurwb.Y2Zypf{animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1)}.edhGSc.u3bW4e>.RpC4Ne>.Bfurwb{animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);transform:scaleX(1)}.edhGSc.FPYHkb>.RpC4Ne{padding-top:24px}.fqp6hd{transform-origin:top left;transform:translate(0,-22px);transition:all .3s cubic-bezier(0.4,0,0.2,1);transition-property:color,top,-webkit-transform;transition-property:color,top,transform;transition-property:color,top,transform,-webkit-transform;color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-size:16px;pointer-events:none;position:absolute;top:100%;width:100%}.edhGSc.u3bW4e>.RpC4Ne>.fqp6hd,.edhGSc.CDELXb>.RpC4Ne>.fqp6hd,.edhGSc.LydCob .fqp6hd{transform:scale(0.75);top:16px}.edhGSc.dm7YTc>.RpC4Ne>.fqp6hd{color:rgba(255,255,255,.38)}.edhGSc.u3bW4e>.RpC4Ne>.fqp6hd,.edhGSc.u3bW4e.dm7YTc>.RpC4Ne>.fqp6hd{color:#4285f4}.F1pOBe{color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;max-width:100%;overflow:hidden;pointer-events:none;position:absolute;bottom:3px;text-overflow:ellipsis;white-space:nowrap}.edhGSc.dm7YTc .F1pOBe{color:rgba(255,255,255,.38)}.edhGSc.CDELXb>.RpC4Ne>.F1pOBe{display:none}.S1BUyf{font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:16px;margin-left:auto;padding-left:16px;padding-top:8px;pointer-events:none;text-align:right;color:rgba(0,0,0,.38);white-space:nowrap}.edhGSc.dm7YTc>.S1BUyf{color:rgba(255,255,255,.38)}.edhGSc.wrxyb{padding-bottom:4px}.v6odTb,.YElZX:not(:empty){-moz-box-flex:1;-moz-box-flex:1 1 auto;flex:1 1 auto;font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;min-height:16px;padding-top:8px}.edhGSc.wrxyb .jE8NUc{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.YElZX{pointer-events:none}.v6odTb{color:#d50000}.edhGSc.dm7YTc .v6odTb{color:#ff6e6e}.YElZX{opacity:.3}.edhGSc.k0tWj .YElZX,.edhGSc:not(.k0tWj) .YElZX:not(:empty)+.v6odTb{display:none}@keyframes quantumWizPaperInputRemoveUnderline{0%{transform:scaleX(1);opacity:1}to{transform:scaleX(1);opacity:0}}@keyframes quantumWizPaperInputAddUnderline{0%{transform:scaleX(0)}to{transform:scaleX(1)}}.LsSwGf{-moz-user-select:none;-moz-box-sizing:content-box;box-sizing:content-box;cursor:pointer;display:inline-block;height:20px;outline:none;position:relative;vertical-align:middle;width:37px;z-index:0}.LsSwGf[aria-disabled=true]{cursor:default}.E7QdY{-moz-transition:border-color .3s ease;transition:border-color .3s ease;border:10px solid #fafafa;-moz-border-radius:100%;border-radius:100%;position:absolute;-moz-box-shadow:0px 1px 3px rgba(0,0,0,.4);box-shadow:0px 1px 3px rgba(0,0,0,.4)}[aria-checked=true] .E7QdY{border-color:#009688}[aria-disabled=true] .E7QdY{border-color:#bdbdbd}.rbsY8b{transition:-webkit-transform .06s ease;transition:transform .06s ease;transition:transform .06s ease,-webkit-transform .06s ease}.LsSwGf.N2RpBe>.rbsY8b{-moz-transform:translate(17px);transform:translate(17px)}.LsSwGf.B6Vhqe>.rbsY8b{-moz-transform:translate(8.5px);transform:translate(8.5px)}.hh4xKf{-moz-transition:border-color .3s ease;transition:border-color .3s ease;border:7px solid #b9b9b9;-moz-border-radius:7px;border-radius:7px;position:absolute;top:3px;width:23px}[aria-checked=true]>.hh4xKf{border-color:rgba(0,150,136,0.502)}[aria-disabled=true]>.hh4xKf{border-color:#b9b9b9}[aria-checked=mixed] .E7QdY{border-color:#f4b400}[aria-checked=mixed] .hh4xKf{border-color:#e0e0e0}[aria-checked=mixed] .YGFwk{left:8.5px}.YGFwk{-moz-transform:scale(2.5);transform:scale(2.5);-moz-transition:opacity 0.15s ease,left 0.3s ease;transition:opacity 0.15s ease,left 0.3s ease;background-color:rgba(0,0,0,0.2);-moz-border-radius:100%;border-radius:100%;height:20px;left:0;opacity:0;outline:.1px solid transparent;pointer-events:none;position:absolute;width:20px;z-index:-1}.qs41qe>.YGFwk{-moz-animation:quantumWizRadialInkSpread .3s;animation:quantumWizRadialInkSpread .3s;animation-fill-mode:forwards;opacity:1}[aria-checked=true]>.YGFwk{left:17px}.i9xfbb>.YGFwk{background-color:rgba(0,150,136,0.2)}.u3bW4e>.YGFwk{-moz-animation:quantumWizRadialInkFocusPulse .7s infinite alternate;animation:quantumWizRadialInkFocusPulse .7s infinite alternate;background-color:rgba(0,150,136,0.2);opacity:1}.Q2P1Eb{-moz-user-select:none;-moz-transition:background-color .1s ease;transition:background-color .1s ease;cursor:pointer;display:block;font-size:14px;font-weight:500;outline:none;overflow:hidden;padding:8px 16px;position:relative}.Q2P1Eb.qs41qe,.Q2P1Eb:focus{background-color:rgba(153,153,153,.2)}.Q2P1Eb.RDPZE{color:rgba(68,68,68,0.502)}.kYtXye .bFjUmb-Ysl7Fe.kRqvHe{background-color:#a1c2fa}.kYtXye .bFjUmb-Wvd9Cc.kRqvHe{background-color:#3b78e7}.eejsDc{overflow-y:auto}.rFrNMe.dm7YTc .cXrdqd{background-color:white}.rFrNMe.dm7YTc:not([disabled]):focus .AxOyFc{color:white}.jBmls .oKubKe{font:0.8125rem "Roboto",Helvetica,Arial,sans-serif;padding-bottom:0.5rem;padding-top:0.5rem}.V6WXSe.CCJ0ld-Jup3Tc{z-index:1192}.c7fp5b{line-height:0}.JRtysb{display:block;height:auto;line-height:0;width:auto}.JRtysb .snByac.snByac{margin:8px}.JRtysb,.mUbCce{flex-shrink:0}.MhXXcc{line-height:0}.fKz7Od,.WzwrXb:not(.K2mXPb){opacity:0.54;transition:opacity 150ms cubic-bezier(0.4,0,0.2,1)}.fKz7Od.RDPZE,.WzwrXb.RDPZE:not(.K2mXPb){opacity:0.26}.fKz7Od:not(.RDPZE):hover,.WzwrXb:not(.RDPZE):not(.K2mXPb):hover{opacity:0.87}.fKz7Od.u3bW4e,.WzwrXb.u3bW4e:not(.K2mXPb),.WzwrXb.iWO5td:not(.K2mXPb){opacity:1}.ZDSs1:not(:hover),.ueScFe:not(:hover),.p9Nwte:not(:hover),.VsxsTb:not(:hover){color:#fff;fill:#fff}.p9Nwte.RDPZE,.ZDSs1.RDPZE{color:#fff;opacity:0.54}.jgvuAb:not(.ybOdnf) .eU809d{border-color:#9e9e9e transparent;border-width:5px 5px 0;top:16px}.jgvuAb.RDPZE .eU809d{border-color:#bdbdbd transparent}.zZhnYe .snByac{margin:0.5rem 1rem}.fKz7Od .TpQm9d{color:black}.p9Nwte .TpQm9d{color:white}.onkcGd,.onkcGd:visited,.etFl5b,.etFl5b:visited,.Vx8Sxd,.Vx8Sxd:visited,.eL9Cfb,.eL9Cfb:visited,.L5mE7d,.L5mE7d:visited,.OGhwGf,.OGhwGf:visited{cursor:pointer;text-decoration:none}.onkcGd,.onkcGd:visited,.OGhwGf,.OGhwGf:visited{color:#333}.FKF6mc{color:#1a73e8}.onkcGd:hover,.onkcGd:focus,.Vx8Sxd:hover,.Vx8Sxd:focus,.etFl5b:hover,.etFl5b:focus,.eL9Cfb:hover,.eL9Cfb:focus,.L5mE7d:hover,.L5mE7d:focus,.OGhwGf:hover,.OGhwGf:focus{outline:none;text-decoration:underline}.onkcGd:hover,.onkcGd:focus,.etFl5b,.etFl5b:visited,.etFl5b:hover,.etFl5b:focus,.eL9Cfb,.eL9Cfb:visited,.eL9Cfb:hover,.eL9Cfb:focus,.L5mE7d,.L5mE7d:visited,.L5mE7d:hover,.L5mE7d:focus,.OGhwGf:hover,.OGhwGf:focus{color:#1a73e8}.Vx8Sxd,.Vx8Sxd:visited,.Vx8Sxd:hover,.Vx8Sxd:focus{color:#fff}.DyGAsf{max-width:21rem}.UtYN2b{max-width:29rem}.SoH8bd{max-width:37rem}.DyGAsf p,.UtYN2b p,.SoH8bd p{margin-bottom:1em}.DyGAsf p:last-child,.UtYN2b p:last-child,.SoH8bd p:last-child{margin-bottom:0}.e8E4Gb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;height:100%}.YVvGBb{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;display:block}.zDK4rb{word-break:break-word}.pco8Kc{display:block;overflow:hidden;overflow-wrap:break-word}.tkmmwb{align-self:flex-start;-moz-border-radius:50%;border-radius:50%;flex-shrink:0;max-height:75px;max-width:75px;vertical-align:middle}.xAhNjc{align-self:center;-moz-border-radius:50%;border-radius:50%;flex-shrink:0;height:2.5rem;margin-right:1rem;vertical-align:middle;width:2.5rem}.j8gm8{visibility:hidden}.L3bAHe{padding:1.5rem}@media (max-width:30em){.L3bAHe{padding:0.5rem}}.G0o5Ac{list-style:disc;padding-left:40px}.FUvKMe{color:rgba(0,0,0,.87)}.OyJCve{color:rgba(0,0,0,.549)}.DPvwYc{font-size:1.5rem;-moz-user-select:none}.DwazCc{font-size:1.125rem}.vUBwW{-moz-border-radius:50%;border-radius:50%;color:rgba(255,255,255,.87);flex-shrink:0;font-size:1rem;height:2rem;line-height:2rem;text-align:center;width:2rem}.vUBwW .DPvwYc{color:white}.oxacD.mUbCce,.oxacD.Y5FYJe,.oxacD.yHy1rc{margin:-12px;display:block}.oxacD.JRtysb,.oxacD.O0WRkf,.oxacD.UQuaGc{display:block;margin:-8px}.oxacD.UQuaGc.cd29Sd{margin:-8px -16px -8px -12px}.oxacD.ksBjEc{margin:-6px -8px -6px -8px}.I2XGyb.jgvuAb{margin-left:-1rem}.tnmqXd{max-width:none}.V1uRod.VfPpkd-MPu53c{margin:-0.25rem 0}@media (max-width:30em){.V1uRod.VfPpkd-MPu53c{margin-left:-0.25rem}}.LBlAUc{margin-bottom:1.5rem}@media (max-width:30em){.LBlAUc{margin-bottom:0.5rem}}.raZwr{margin-bottom:2rem}@media (max-width:30em){.raZwr{margin-bottom:1.5rem}}.QRiHXd{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row}.ZFZEWb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center}.bxp7vf{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center}.vgYYId{box-sizing:border-box;height:100%;width:100%}.Vv9Gs{-moz-box-flex:1 0 2rem;flex:1 0 2rem}.iXypXd{-moz-box-flex:1 0 1.5rem;flex:1 0 1.5rem}.Nmpzvc{-moz-box-flex:1 0 1rem;flex:1 0 1rem}.fPqOAb{-moz-box-flex:1 0 0.5rem;flex:1 0 0.5rem}img[src='']{visibility:hidden}.WG5SSb{max-height:0.0625rem;max-width:0.0625rem;opacity:.001;pointer-events:none;position:absolute;visibility:visible}.PazDv{font-size:0.0625rem;height:0.0625rem;line-height:1;opacity:.001;overflow:hidden;position:absolute;width:0.0625rem}@keyframes hrFadeIn{0%{opacity:0}to{opacity:1}}@keyframes hrRippleTransform{0%{transform:scale(0)}to{transform:scale(1)}}.ULzZ3{-moz-border-radius:50%;border-radius:50%;bottom:-100%;height:300%;left:-100%;opacity:0;position:absolute;top:-100%;right:-100%;width:300%}.FAtkpf{align-items:center;height:-moz-calc(100vh - 4rem);height:calc(100vh - 4rem);display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-flow:column;justify-content:center;left:0;position:absolute;right:0;top:4rem}.FAtkpf>*{flex-shrink:0}em,strong{font-weight:500;font-style:normal}.rwnykc{color:rgba(0,0,0,.549);font-size:2.8125rem;font-weight:400;line-height:3rem}.nk37z{color:rgba(0,0,0,.87);font-size:1.25rem;font-weight:500;line-height:1.75rem}.CHXfbe{color:rgba(0,0,0,.549);font-size:1.25rem;font-weight:500;line-height:1.75rem}.udxSmc{color:rgba(0,0,0,.549);font-size:0.75rem;font-weight:400}.i9glDf{color:rgba(0,0,0,.87);font-size:0.9375rem;font-weight:500}.VIwAmc{color:rgba(0,0,0,.549);font-size:0.9375rem;font-weight:400}.Evt7cb,.Evt7cb:visited{color:rgba(0,0,0,.87);font-size:0.8125rem;font-weight:500;line-height:1.5rem}.KATzH,.KATzH:visited{color:rgba(0,0,0,.549);font-size:0.8125rem;font-weight:500;line-height:1.5rem}.lziZub,.lziZub:visited{color:rgba(0,0,0,.87);font-size:0.8125rem;font-weight:400;line-height:1.25rem}.IMvYId,.IMvYId:visited{color:rgba(0,0,0,.549);font-size:0.8125rem;font-weight:400;line-height:1.25rem}@media (max-width:40em){.s7bwNb,.i9glDf,.VIwAmc{font-size:1rem}.udxSmc,.DWxSed,.x4sAde,.EWXgRe,.Evt7cb,.KATzH,.lziZub,.IMvYId,.vHZOhb{font-size:0.875rem}}.vzcr8{color:#2e7d32}.Kma9Mb{color:#d50000}.neggzd{color:transparent;cursor:default;text-shadow:0 0 .7em rgba(0,0,0,.549);-moz-user-select:none}iframe[name="google-hats-survey"]{z-index:9998}.iph-dialog-content ul{list-style:disc;margin:1em 0;padding-left:1.5rem}.iph-dialog-content a[href]:focus{background-color:rgba(0,0,0,.1);border-radius:0.125rem;margin:-0.25rem -0.5rem;padding:0.25rem 0.5rem}.a5kY4d{border:0.0625rem solid #e0e0e0;-moz-border-radius:1.1875rem;border-radius:1.1875rem;box-flex:1;flex-grow:1;-moz-flex-wrap:wrap;flex-wrap:wrap;justify-content:flex-end;margin:0.0625rem}.a5kY4d:focus-within{border-width:0.125rem;margin:0}.nxIm7c{box-flex:1;flex-grow:1;overflow:hidden;padding:0.375rem 0.9375rem}.vaUyHb{font-family:"Google Sans Display",Roboto,Arial,sans-serif;font-size:2.75rem;font-weight:400;line-height:3.25rem}@media (max-width:40em){.vaUyHb{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:2.25rem;font-weight:400;line-height:2.75rem}}.YrFhrf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:2.25rem;font-weight:400;line-height:2.75rem;color:#3c4043}.YrFhrf-ZoZQ1{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:2.25rem;font-weight:500;line-height:2.75rem;color:#fff}@media (max-width:40em){.YrFhrf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.75rem;font-weight:400;line-height:2.25rem}.YrFhrf-ZoZQ1{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.75rem;font-weight:500;line-height:2.25rem}}.B7SYid{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:2rem;font-weight:400;line-height:2.5rem}@media (max-width:40em){.B7SYid{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.75rem;font-weight:400;line-height:2.25rem}}.kGNarb{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.75rem;font-weight:400;line-height:2.25rem}.BYh5cb{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.5rem;font-weight:400;line-height:2rem}.z3vRcc-ZoZQ1{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;line-height:1.75rem;color:#fff}.z3vRcc{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;line-height:1.75rem;color:#3c4043}.z3vRcc-J3yWx{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;line-height:1.75rem;color:#5f6368}@media (max-width:40em){.z3vRcc-ZoZQ1,.z3vRcc,.z3vRcc-J3yWx{letter-spacing:.00625em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1rem;font-weight:400;line-height:1.5rem}}.WOPwXe{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.125rem;font-weight:400;line-height:1.5rem;color:#3c4043}.WOPwXe-Wvd9Cc{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.125rem;font-weight:500;line-height:1.5rem;color:#3c4043}.A6dC2c{letter-spacing:.00625em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1rem;font-weight:500;line-height:1.5rem;color:#3c4043}.EZrbnd{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#3c4043;text-transform:none}.asQXV{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#3c4043}.iLjzDc{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#5f6368}.asQXV-FGzYL{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:400;line-height:1.25rem;color:#3c4043}.lYU7F{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#c5221f}.EhRlC{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#1e8e3e}.gJk24c{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#1967d2}.pO05gd{letter-spacing:.00625em;font-family:Roboto,Arial,sans-serif;font-size:1rem;font-weight:400;line-height:1.5rem;color:#3c4043}.tLDEHd{letter-spacing:.01428571em;font-family:Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:400;line-height:1.25rem;color:#3c4043}.tLDEHd-Wvd9Cc{letter-spacing:.01428571em;font-family:Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#5f6368}.cSyPgb{letter-spacing:.01428571em;font-family:Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:400;line-height:1.25rem;color:#5f6368}.dDKhVc{letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:0.75rem;font-weight:400;line-height:1rem;color:#5f6368}.dDKhVc-Wvd9Cc{letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:0.75rem;font-weight:500;line-height:1rem;color:#5f6368}.T8rTjd{letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:0.75rem;font-weight:400;line-height:1rem;color:#5f6368;display:inline-block}.M1rIWd{letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:0.75rem;font-weight:400;line-height:1rem;color:#b31412}.ViCi4{letter-spacing:.01785714em;font-family:Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;color:#3c4043}.Aopndd{background-color:#fff;border:0.0625rem solid #dadce0;-moz-border-radius:0.5rem;border-radius:0.5rem;overflow:hidden}.GWZ7yf{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);border-radius:0.5rem;overflow:hidden}.n0p5v{padding:1.5rem}@media (max-width:30em){.n0p5v{padding:0.5rem}}.xSP5ic,.xSP5ic.yHy1rc{color:#5f6368;fill:#5f6368}.e0pgvc,.xSP5ic.e0pgvc{color:#9aa0a6;fill:#9aa0a6}.uwbd3d svg{width:1.125rem;height:1.125rem}.m1PbN{color:#fff;fill:#fff}.yJ0xsb.UQuaGc:not(.RDPZE) .TpQm9d{background:none}.LKmtKf:hover,.S6Vdac:hover{background-color:rgba(32,33,36,0.039)}.CAntkd:focus,.S6Vdac:focus{background-color:rgba(32,33,36,0.122)}.S3R4yc .snByac{fill:currentcolor}.tUJKGd:not(:first-child){border-top:0.0625rem solid #e0e0e0}.tUJKGd:hover,.tUJKGd:focus-within{-moz-border-radius:0.5rem;border-radius:0.5rem;overflow:hidden}.tUJKGd:not(:first-child):hover,.tUJKGd:not(:first-child):focus-within,.tUJKGd:hover+.tUJKGd,.tUJKGd:focus-within+.tUJKGd{border-top-color:transparent}.uO32ac{height:4.5rem}.iph-dialog.iph-dialog{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);border-radius:0.5rem;overflow:hidden}.iph-dialog .iph-dialog-title{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;line-height:1.75rem}.iph-dialog.iph-dialog button{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;text-transform:none}.cLpBac{background:#f8f9fa;padding:12px 0}.cLpBac .Fxmcue{padding-left:1rem}.cLpBac.TuHiFd .snByac,.cLpBac.REtOWc .snByac{width:100%}.QTD2uf{border:0.0625rem solid #dadce0;-moz-border-radius:0.5rem;border-radius:0.5rem;display:block;width:100%}.QTD2uf .OA0qNb{max-width:100%}.QTD2uf.QTD2uf .oJeWuf{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;display:block}.TNy2be.TNy2be.TNy2be{margin-bottom:0.4375rem;margin-right:0.875rem}.dkNZte{background:#e8eaed;-moz-border-radius:0.25rem;border-radius:0.25rem;line-height:1.5rem;margin-left:1rem;padding:0 0.5rem}.oQOrod{margin:0 0.25rem}.zg38Fd{display:inline-block;margin-left:0.5rem;vertical-align:sub}.slQh3d{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin:1rem 0}.Yxrrpd{margin-right:0.5rem}.EmVfjc{display:inline-block;position:relative;width:28px;height:28px}.Cg7hO{position:absolute;width:0;height:0;overflow:hidden}.xu46lf{width:100%;height:100%}.EmVfjc.qs41qe .xu46lf{animation:spinner-container-rotate 1568ms linear infinite}.ir3uv{position:absolute;width:100%;height:100%;opacity:0}.uWlRce{border-color:#4285f4}.GFoASc{border-color:#db4437}.WpeOqd{border-color:#f4b400}.rHV3jf{border-color:#0f9d58}.EmVfjc.qs41qe .ir3uv.uWlRce{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-blue-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.EmVfjc.qs41qe .ir3uv.GFoASc{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-red-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.EmVfjc.qs41qe .ir3uv.WpeOqd{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-yellow-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.EmVfjc.qs41qe .ir3uv.rHV3jf{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-green-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.HBnAAc{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;top:0;left:45%;width:10%;height:100%;overflow:hidden;border-color:inherit}.HBnAAc .X6jHbb{width:1000%;left:-450%}.xq3j6{display:inline-block;position:relative;width:50%;height:100%;overflow:hidden;border-color:inherit}.xq3j6 .X6jHbb{width:200%}.X6jHbb{position:absolute;top:0;right:0;bottom:0;left:0;-moz-box-sizing:border-box;box-sizing:border-box;height:100%;border-width:3px;border-style:solid;border-color:inherit;border-bottom-color:transparent;-moz-border-radius:50%;border-radius:50%;animation:none}.xq3j6.ERcjC .X6jHbb{border-right-color:transparent;transform:rotate(129deg)}.xq3j6.dj3yTd .X6jHbb{left:-100%;border-left-color:transparent;transform:rotate(-129deg)}.EmVfjc.qs41qe .xq3j6.ERcjC .X6jHbb{animation:spinner-left-spin 1333ms cubic-bezier(0.4,0,0.2,1) infinite both}.EmVfjc.qs41qe .xq3j6.dj3yTd .X6jHbb{animation:spinner-right-spin 1333ms cubic-bezier(0.4,0,0.2,1) infinite both}.EmVfjc.sf4e6b .xu46lf{animation:spinner-container-rotate 1568ms linear infinite,spinner-fade-out 400ms cubic-bezier(0.4,0,0.2,1)}@keyframes spinner-container-rotate{to{transform:rotate(360deg)}}@keyframes spinner-fill-unfill-rotate{12.5%{transform:rotate(135deg)}25%{transform:rotate(270deg)}37.5%{transform:rotate(405deg)}50%{transform:rotate(540deg)}62.5%{transform:rotate(675deg)}75%{transform:rotate(810deg)}87.5%{transform:rotate(945deg)}to{transform:rotate(1080deg)}}@keyframes spinner-blue-fade-in-out{0%{opacity:.99}25%{opacity:.99}26%{opacity:0}89%{opacity:0}90%{opacity:.99}to{opacity:.99}}@keyframes spinner-red-fade-in-out{0%{opacity:0}15%{opacity:0}25%{opacity:.99}50%{opacity:.99}51%{opacity:0}}@keyframes spinner-yellow-fade-in-out{0%{opacity:0}40%{opacity:0}50%{opacity:.99}75%{opacity:.99}76%{opacity:0}}@keyframes spinner-green-fade-in-out{0%{opacity:0}65%{opacity:0}75%{opacity:.99}90%{opacity:.99}to{opacity:0}}@keyframes spinner-left-spin{0%{transform:rotate(130deg)}50%{transform:rotate(-5deg)}to{transform:rotate(130deg)}}@keyframes spinner-right-spin{0%{transform:rotate(-130deg)}50%{transform:rotate(5deg)}to{transform:rotate(-130deg)}}@keyframes spinner-fade-out{0%{opacity:.99}to{opacity:0}}.f0kHoc{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;justify-content:center;width:100%}.aP3ZPb{height:0.25rem;overflow:hidden;position:relative;width:100%}.bNpzdf{animation:hrLoadingIndicatorMove 1400ms infinite,hrLoadingIndicatorVaryWidth 1300ms infinite;animation-timing-function:cubic-bezier(0.4,0.0,0.2,1);transform-origin:right top;left:-60%;position:absolute}.G1kKid{animation:hrLoadingIndicatorMove 1400ms infinite cubic-bezier(0.4,0.0,0.2,1);animation-delay:700ms;left:-60%;position:absolute;width:60%}.Po14Kd{background-color:#fff}.BWOvob{background-color:#a0c1fc}@keyframes hrLoadingIndicatorMove{0%{left:-60%}to{left:100%}}@keyframes hrLoadingIndicatorVaryWidth{0%{width:60%}10%{width:60%}66%{width:1%}to{width:60%}}.IrxBzb,.IrxBzb:focus,.IrxBzb:visited{color:inherit;display:block;fill:inherit;outline:none;stroke:inherit;text-decoration:none}.uArJ5e.u3bW4e{outline:1px solid transparent}.NMm5M{fill:currentColor;flex-shrink:0}html[dir=rtl] .hhikbc{transform:scaleX(-1)}.j70YMc ol,.j70YMc ul{margin:1em 0;padding-left:40px}.j70YMc ol{list-style:decimal}.j70YMc ul{list-style:disc}.q1Kmyc{border:.0625rem solid rgb(218,220,224);border-radius:1.5rem;-moz-box-flex:1;flex-grow:1;flex-wrap:wrap;-moz-box-pack:end;justify-content:flex-end;margin:.0625rem}.q1Kmyc:focus-within{border-width:.125rem;margin:0}.pPgY8b:not(:focus-within) .CIy9F{display:none}.pPgY8b:not(:focus-within) .snByac{top:.625rem}.pPgY8b:not(:focus-within) .I9OJHe{padding:.375rem 1rem}.pPgY8b .snByac{font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400;color:rgb(128,134,139)}.pPgY8b .CIy9F{border-radius:0 0 1rem 1rem;padding-left:.5rem}.pPgY8b .mIZh1c,.pPgY8b .cXrdqd{display:none}.xVPuB .I9OJHe,.vnnr5e .I9OJHe{-moz-border-radius:4px 4px 0 0;border-radius:4px 4px 0 0;padding:10px 16px}.xVPuB .I9OJHe.vTcY1d,.vnnr5e .I9OJHe.vTcY1d{padding-top:22px}.xVPuB.RDPZE .I9OJHe,.vnnr5e.RDPZE .I9OJHe{background-color:rgba(248,249,250,.38)}.xVPuB .snByac,.vnnr5e .snByac{color:#5f6368;padding-left:16px;top:18px}.vnnr5e.u3bW4e .I9OJHe.vTcY1d .snByac,.vnnr5e.CDELXb .I9OJHe.vTcY1d .snByac{transform:scale(0.75) translateX(5px) translateY(-27px)}.xVPuB .KRoqRc,.vnnr5e .KRoqRc{margin-top:2px}.xVPuB .mIZh1c,.vnnr5e .mIZh1c{background-color:#80868b}.xVPuB .mIZh1c,.xVPuB .cXrdqd,.vnnr5e .mIZh1c,.vnnr5e .cXrdqd{bottom:-41px}.xVPuB.u3bW4e .snByac{font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400;top:12px}.vnnr5e .I9OJHe,.vnnr5e .CIy9F{background-color:#f8f9fa}.vnnr5e:not(.RDPZE):hover .I9OJHe,.vnnr5e:not(.RDPZE):hover .CIy9F{background-color:#f1f3f4}.xVPuB .Aworge,.vnnr5e .Aworge{color:#5f6368;height:34px;opacity:1;width:36px}.zuzKle.xVPuB,.zuzKle.vnnr5e{width:100%}.a5lbif{height:2rem;width:2rem;margin-right:1rem}.YfRA6b{align-self:start;padding:.375rem 0}.AI7uec{align-self:auto}.RFmjW{max-width:calc(100% - 2.75rem)}.GngEL{max-width:calc(100% - 5.75rem)}.yUZA2d{max-width:calc(100% - 3rem)}.apsLYe{align-self:flex-end;margin-right:.25rem}.C83nhf{padding-bottom:.25rem}.T8tcPb{height:2.25rem;width:2.25rem}.T8tcPb .GmuOkf{left:.125rem}.apsLYe.apsLYe .f0kHoc{margin:.25rem .5rem .5rem .25rem}.apsLYe .EmVfjc{height:1.125rem;margin:mult(sub(SAVE_BUTTON_SIZE,1.125rem),.5);width:1.125rem}body{color:rgba(0,0,0,.87);font-family:"Roboto",Helvetica,Arial,sans-serif;font-size:0.8125rem;font-weight:400;line-height:1.25rem;margin:0;min-width:18.75rem}@media (max-width:40em){body{font-size:0.875rem}}h1,h2,h3,h4,h5,h6{font-size:inherit;font-weight:inherit;margin:0}input,textarea,keygen,select,button{font:inherit}:focus{outline:1px solid transparent}ul,ol{list-style:none;margin:0;padding:0}p{margin:0}.kFwPee{height:100%}.ydMMEb{width:100%}.SSPGKf{display:block;overflow-y:hidden;z-index:1}.eejsDc{overflow-y:auto}.MCcOAc{bottom:0;left:0;position:absolute;right:0;top:0;overflow:hidden;z-index:1}.MCcOAc>.pGxpHc{flex-shrink:0;box-flex:0;flex-grow:0}.IqBfM>.HLlAHb{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:60px;position:absolute;right:16px;top:0;z-index:9999}.VUoKZ{display:none;position:absolute;top:0;left:0;right:0;height:3px;z-index:1001}.TRHLAc{position:absolute;top:0;left:0;width:25%;height:100%;background:#68e;transform:scaleX(0);transform-origin:0 0}.mIM26c .VUoKZ{display:block}.mIM26c .TRHLAc{animation:boqChromeapiPageProgressAnimation 1s infinite;animation-timing-function:cubic-bezier(0.4,0.0,1,1);animation-delay:.1s}.ghyPEc .VUoKZ{position:fixed}@keyframes boqChromeapiPageProgressAnimation{0%{transform:scaleX(0)}50%{transform:scaleX(5)}to{transform:scaleX(5) translateX(100%)}}c-wiz{contain:style}c-wiz>c-data{display:none}c-wiz.rETSD{contain:none}c-wiz.Ubi8Z{contain:layout style}.Qks78e{overflow:hidden}.JtDYBc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-shrink:0;justify-content:center;margin-right:1.5rem;width:2rem}.TGnLfc{color:#fff;line-height:2rem;text-transform:uppercase}.HbHNgd{overflow:hidden}.VfPpkd-I9GLp-yrriRe{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit);color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87));display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center;vertical-align:middle}.VfPpkd-I9GLp-yrriRe[hidden]{display:none}.VfPpkd-I9GLp-yrriRe>label{margin-left:0;margin-right:auto;padding-left:4px;padding-right:0;-moz-box-ordinal-group:1;order:0}[dir=rtl] .VfPpkd-I9GLp-yrriRe>label,.VfPpkd-I9GLp-yrriRe>label[dir=rtl]{margin-left:auto;margin-right:0}[dir=rtl] .VfPpkd-I9GLp-yrriRe>label,.VfPpkd-I9GLp-yrriRe>label[dir=rtl]{padding-left:0;padding-right:4px}.VfPpkd-I9GLp-yrriRe-OWXEXe-WrakWd>label{text-overflow:ellipsis;overflow:hidden;white-space:nowrap}.VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d>label{margin-left:auto;margin-right:0;padding-left:0;padding-right:4px;-moz-box-ordinal-group:0;order:-1}[dir=rtl] .VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d>label,.VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d>label[dir=rtl]{margin-left:0;margin-right:auto}[dir=rtl] .VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d>label,.VfPpkd-I9GLp-yrriRe-OWXEXe-fW01td-CpWD9d>label[dir=rtl]{padding-left:4px;padding-right:0}.VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL{-moz-box-pack:justify;justify-content:space-between}.VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL>label{margin:0}[dir=rtl] .VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL>label,.VfPpkd-I9GLp-yrriRe-OWXEXe-fozPsf-t6UvL>label[dir=rtl]{margin:0}.MlG5Jc{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400}.MlG5Jc gm-checkbox[disabled]~.VfPpkd-V67aGc,.MlG5Jc gm-radio[disabled]~.VfPpkd-V67aGc,.MlG5Jc .VfPpkd-MPu53c-OWXEXe-OWB6Me~.VfPpkd-V67aGc,.MlG5Jc .VfPpkd-GCYh9b-OWXEXe-OWB6Me~.VfPpkd-V67aGc{color:rgb(95,99,104)}html[dir=rtl] .giSqbe{transform:scaleX(-1)}@keyframes hrUiDrawerIn{0%{transform:translateX(-19.25rem)}100%{transform:translateX(0)}}@keyframes hrUiDrawerOut{0%{transform:translateX(0)}100%{transform:translateX(-19.25rem)}}@keyframes hrRtlUiDrawerIn{0%{transform:translateX(19.25rem)}100%{transform:translateX(0)}}@keyframes hrRtlUiDrawerOut{0%{transform:translateX(0)}100%{transform:translateX(19.25rem)}}@keyframes hrUiDrawerItemRipple{0%{transform:scale(0)}100%{transform:scale(1)}}.AxPfNe{bottom:0;height:100vh;left:0;opacity:0;overflow:hidden;position:fixed;right:0;top:0;width:100vw;z-index:990}.dgqqXe .AxPfNe,.OMVS8d .AxPfNe{display:none}.ETRkCe{box-shadow:0 4px 4px 0 rgba(60,64,67,.3),0 8px 12px 6px rgba(60,64,67,.15);background-color:#fff;bottom:0;height:100vh;left:0;position:fixed;top:0;width:19rem;z-index:990}.CBSF1e .ETRkCe{transform:translateX(0)}.dgqqXe .ETRkCe{display:none;visibility:hidden}.X1rxSc .ETRkCe{animation:hrUiDrawerIn .3s cubic-bezier(0,0,.2,1) forwards}.OMVS8d .ETRkCe{animation:hrUiDrawerOut .3s cubic-bezier(0,0,.2,1) forwards}[dir=rtl] .X1rxSc .ETRkCe{animation:hrRtlUiDrawerIn .3s cubic-bezier(0,0,.2,1) forwards}[dir=rtl] .OMVS8d .ETRkCe{animation:hrRtlUiDrawerOut .3s cubic-bezier(0,0,.2,1) forwards}.Tabkde{-moz-box-flex:1;flex:1 1 auto;position:relative;width:19rem}.Tabkde:before{background-color:#fff;bottom:0;content:"";left:0;position:absolute;right:0;top:0;z-index:-2}.ideBx{width:19rem;-moz-box-flex:0;flex:0 0 19rem}.Hlw1k .ideBx{display:none}@media (max-width:65.125rem){.ideBx{display:none}}.Du1LZe{height:100%;min-height:0}.OX4Vcb{-moz-box-sizing:border-box;box-sizing:border-box;height:100%;overflow-x:hidden;overflow-y:auto;padding-bottom:.5rem;padding-top:.5rem;width:100%}.Xi8cpb{-moz-box-align:center;align-items:center;cursor:pointer;display:-moz-box;display:flex;height:3.5rem;padding-left:1rem;padding-right:1rem;position:relative}.x2LcDe a.Xi8cpb{text-decoration:none}.Xi8cpb.vG1fDb{height:4rem}.LlcfK{border-radius:0 2rem 2rem 0;bottom:0;left:0;overflow:hidden;position:absolute;right:.5rem;top:0;z-index:-1}.p1KYTc{border-radius:50%;bottom:0;height:300%;left:-100%;position:absolute;top:-100%;right:0;width:300%}.kYtXye .Xi8cpb.qs41qe .LlcfK{background-color:rgba(26,115,232,.12)}.Xi8cpb:hover .LlcfK{background-color:rgba(32,33,36,.04)}.Xi8cpb:focus .LlcfK{background-color:rgba(32,33,36,.08)}.Xi8cpb:active .p1KYTc{animation:hrUiDrawerItemRipple .2s cubic-bezier(0,0,.2,1) forwards;background-color:rgba(26,115,232,.06)}.pkktJb{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;height:2.5rem;padding-left:1rem;padding-right:1rem}.yXVLvd,.JDxyrc{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-flex:0;flex:0 0 auto;-moz-box-pack:center;justify-content:center;width:2.5rem}.oOEg5c{background:rgb(206,234,214);border-radius:52px;color:rgb(13,101,45);font-weight:500;line-height:20px;margin-left:16px;padding:0 6px;text-align:center}.kXvNXe{margin-left:1rem;overflow:hidden}.utCGpd{display:-moz-box;display:flex}.mzwNCf{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;height:4rem;-moz-box-pack:center;justify-content:center}.yCa5be{list-style:none;margin:.5rem 0}.IqJTee{color:#5f6368;font-family:"Product Sans",Arial,Helvetica,sans-serif;font-size:1.38125rem;position:relative;top:-.375rem;text-rendering:optimizeLegibility;-moz-osx-font-smoothing:grayscale}.VfPpkd-JGcpL-uI4vCe-LkdAo,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#6200ee;stroke:var(--mdc-theme-primary,#6200ee)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-JGcpL-uI4vCe-LkdAo,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.VfPpkd-JGcpL-uI4vCe-u014N{stroke:transparent}@keyframes mdc-circular-progress-container-rotate{to{transform:rotate(1turn)}}@keyframes mdc-circular-progress-spinner-layer-rotate{12.5%{transform:rotate(135deg)}25%{transform:rotate(270deg)}37.5%{transform:rotate(405deg)}50%{transform:rotate(540deg)}62.5%{transform:rotate(675deg)}75%{transform:rotate(810deg)}87.5%{transform:rotate(945deg)}100%{transform:rotate(3turn)}}@keyframes mdc-circular-progress-color-1-fade-in-out{from{opacity:.99}25%{opacity:.99}26%{opacity:0}89%{opacity:0}90%{opacity:.99}to{opacity:.99}}@keyframes mdc-circular-progress-color-2-fade-in-out{from{opacity:0}15%{opacity:0}25%{opacity:.99}50%{opacity:.99}51%{opacity:0}to{opacity:0}}@keyframes mdc-circular-progress-color-3-fade-in-out{from{opacity:0}40%{opacity:0}50%{opacity:.99}75%{opacity:.99}76%{opacity:0}to{opacity:0}}@keyframes mdc-circular-progress-color-4-fade-in-out{from{opacity:0}65%{opacity:0}75%{opacity:.99}90%{opacity:.99}to{opacity:0}}@keyframes mdc-circular-progress-left-spin{from{transform:rotate(265deg)}50%{transform:rotate(130deg)}to{transform:rotate(265deg)}}@keyframes mdc-circular-progress-right-spin{from{transform:rotate(-265deg)}50%{transform:rotate(-130deg)}to{transform:rotate(-265deg)}}.VfPpkd-JGcpL-P1ekSe{display:-moz-inline-box;display:inline-flex;position:relative;direction:ltr;line-height:0;transition:opacity .25s 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-JGcpL-uI4vCe-haAclf,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G,.VfPpkd-JGcpL-IdXvz-haAclf,.VfPpkd-JGcpL-QYI5B-pbTTYe{position:absolute;width:100%;height:100%}.VfPpkd-JGcpL-uI4vCe-haAclf{transform:rotate(-90deg)}.VfPpkd-JGcpL-IdXvz-haAclf{font-size:0;letter-spacing:0;white-space:nowrap;opacity:0}.VfPpkd-JGcpL-uI4vCe-LkdAo-Bd00G,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{fill:transparent}.VfPpkd-JGcpL-uI4vCe-LkdAo{transition:stroke-dashoffset .5s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-JGcpL-OcUoKf-TpMipd{position:absolute;top:0;left:47.5%;-moz-box-sizing:border-box;box-sizing:border-box;width:5%;height:100%;overflow:hidden}.VfPpkd-JGcpL-OcUoKf-TpMipd .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{left:-900%;width:2000%;transform:rotate(180deg)}.VfPpkd-JGcpL-lLvYUc-e9ayKc{display:-moz-inline-box;display:inline-flex;position:relative;width:50%;height:100%;overflow:hidden}.VfPpkd-JGcpL-lLvYUc-e9ayKc .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{width:200%}.VfPpkd-JGcpL-lLvYUc-qwU8Me .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{left:-100%}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-uI4vCe-haAclf{opacity:0}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-IdXvz-haAclf{opacity:1}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-IdXvz-haAclf{animation:mdc-circular-progress-container-rotate 1.5682352941176s linear infinite}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-QYI5B-pbTTYe{animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-R6PoUb{animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-1-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-ibL1re{animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-2-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-c5RTEf{animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-3-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-II5mzb{animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-4-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-lLvYUc-LK5yu .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{animation:mdc-circular-progress-left-spin 1333ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-lLvYUc-qwU8Me .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{animation:mdc-circular-progress-right-spin 1333ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-xTMeO{opacity:0}.DU29of{position:relative}.DU29of .VfPpkd-JGcpL-uI4vCe-LkdAo,.DU29of .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#4285f4}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-uI4vCe-LkdAo,.DU29of .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#4285f4}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#ea4335}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#fbbc04}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#34a853}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Mr8B3-V67aGc{height:100%;width:100%;position:absolute;opacity:0;overflow:hidden;z-index:-1}.NZp2ef{background-color:#e8eaed}.VfPpkd-z59Tgd{border-radius:4px;border-radius:var(--mdc-shape-small,4px)}.VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.VfPpkd-Djsh7e-XxIAqe-cGMI2b{border-radius:4px;border-radius:var(--mdc-shape-small,4px)}.VfPpkd-z59Tgd{color:white;color:var(--mdc-theme-text-primary-on-dark,white)}.VfPpkd-z59Tgd{background-color:rgba(0,0,0,.6)}.VfPpkd-MlC99b{color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-light,rgba(0,0,0,.87))}.VfPpkd-IqDDtd{color:rgba(0,0,0,.6)}.VfPpkd-IqDDtd-hSRGPd{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{background-color:#fff}.VfPpkd-z59Tgd{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit)}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{box-shadow:0 3px 1px -2px rgba(0,0,0,.2),0 2px 2px 0 rgba(0,0,0,.14),0 1px 5px 0 rgba(0,0,0,.12);border-radius:4px;line-height:20px}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-z59Tgd .VfPpkd-MlC99b{display:block;margin-top:0;line-height:20px;-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-subtitle2-font-size,.875rem);line-height:1.375rem;line-height:var(--mdc-typography-subtitle2-line-height,1.375rem);font-weight:500;font-weight:var(--mdc-typography-subtitle2-font-weight,500);letter-spacing:.0071428571em;letter-spacing:var(--mdc-typography-subtitle2-letter-spacing,.0071428571em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle2-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle2-text-transform,inherit)}.VfPpkd-z59Tgd .VfPpkd-MlC99b::before{display:inline-block;width:0;height:24px;content:"";vertical-align:0}.VfPpkd-z59Tgd .VfPpkd-IqDDtd{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit)}.VfPpkd-z59Tgd{word-break:break-all;word-break:var(--mdc-tooltip-word-break,normal);overflow-wrap:anywhere}.VfPpkd-suEOdc-OWXEXe-eo9XGd-RCfa3e .VfPpkd-z59Tgd-OiiCO{transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),transform .15s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-suEOdc-OWXEXe-ZYIfFd-RCfa3e .VfPpkd-z59Tgd-OiiCO{transition:opacity 75ms 0ms cubic-bezier(.4,0,1,1)}.VfPpkd-suEOdc{position:fixed;display:none;z-index:9}.VfPpkd-suEOdc-sM5MNb-OWXEXe-nzrxxc{position:relative}.VfPpkd-suEOdc-OWXEXe-TSZdd,.VfPpkd-suEOdc-OWXEXe-eo9XGd,.VfPpkd-suEOdc-OWXEXe-ZYIfFd{display:-moz-inline-box;display:inline-flex}.VfPpkd-suEOdc-OWXEXe-TSZdd.VfPpkd-suEOdc-OWXEXe-nzrxxc,.VfPpkd-suEOdc-OWXEXe-eo9XGd.VfPpkd-suEOdc-OWXEXe-nzrxxc,.VfPpkd-suEOdc-OWXEXe-ZYIfFd.VfPpkd-suEOdc-OWXEXe-nzrxxc{display:inline-block;left:-320px;position:absolute}.VfPpkd-z59Tgd{line-height:16px;padding:4px 8px;min-width:40px;max-width:200px;min-height:24px;max-height:40vh;-moz-box-sizing:border-box;box-sizing:border-box;overflow:hidden;text-align:center}.VfPpkd-z59Tgd::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-z59Tgd::before{border-color:CanvasText}}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{-moz-box-align:start;align-items:flex-start;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;min-height:24px;min-width:40px;max-width:320px;position:relative}.VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd{text-align:left}[dir=rtl] .VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd,.VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd[dir=rtl]{text-align:right}.VfPpkd-z59Tgd .VfPpkd-MlC99b{margin:0 8px}.VfPpkd-z59Tgd .VfPpkd-IqDDtd{max-width:184px;margin:8px;text-align:left}[dir=rtl] .VfPpkd-z59Tgd .VfPpkd-IqDDtd,.VfPpkd-z59Tgd .VfPpkd-IqDDtd[dir=rtl]{text-align:right}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd .VfPpkd-IqDDtd{max-width:304px;align-self:stretch}.VfPpkd-z59Tgd .VfPpkd-IqDDtd-hSRGPd{text-decoration:none}.VfPpkd-suEOdc-OWXEXe-nzrxxc-LQLjdd,.VfPpkd-IqDDtd,.VfPpkd-MlC99b{z-index:1}.VfPpkd-z59Tgd-OiiCO{opacity:0;transform:scale(.8);will-change:transform,opacity}.VfPpkd-suEOdc-OWXEXe-TSZdd .VfPpkd-z59Tgd-OiiCO{transform:scale(1);opacity:1}.VfPpkd-suEOdc-OWXEXe-ZYIfFd .VfPpkd-z59Tgd-OiiCO{transform:scale(1)}.VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.VfPpkd-Djsh7e-XxIAqe-cGMI2b{position:absolute;height:24px;width:24px;transform:rotate(35deg) skewY(20deg) scaleX(.9396926208)}.VfPpkd-Djsh7e-XxIAqe-ma6Yeb .VfPpkd-BFbNVe-bF1uUb,.VfPpkd-Djsh7e-XxIAqe-cGMI2b .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-Djsh7e-XxIAqe-cGMI2b{box-shadow:0 3px 1px -2px rgba(0,0,0,.2),0 2px 2px 0 rgba(0,0,0,.14),0 1px 5px 0 rgba(0,0,0,.12);outline:1px solid transparent;z-index:-1}@media screen and (forced-colors:active){.VfPpkd-Djsh7e-XxIAqe-cGMI2b{outline-color:CanvasText}}.EY8ABd{z-index:2101}.EY8ABd .VfPpkd-z59Tgd{background-color:#3c4043;color:#e8eaed}.EY8ABd .VfPpkd-MlC99b,.EY8ABd .VfPpkd-IqDDtd{color:#3c4043}.EY8ABd .VfPpkd-IqDDtd-hSRGPd{color:#1a73e8}.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{background-color:#fff}.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-MlC99b{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{-moz-border-radius:8px;border-radius:8px}.ziykHb{z-index:2101}.ziykHb .VfPpkd-z59Tgd{background-color:#3c4043;color:#e8eaed}.ziykHb .VfPpkd-MlC99b,.ziykHb .VfPpkd-IqDDtd{color:#3c4043}.ziykHb .VfPpkd-IqDDtd-hSRGPd{color:#1a73e8}.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{background-color:#fff}.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-MlC99b{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{-moz-border-radius:8px;border-radius:8px}.EY8ABd-OWXEXe-TAWMXe{position:absolute;left:-10000px;top:auto;width:1px;height:1px;overflow:hidden;-moz-user-select:none;-moz-user-select:none}.ZSrdFd{-moz-user-select:none;cursor:pointer;display:inline-block;text-decoration:none}.ZSrdFd:focus{outline:none}.ZSrdFd:hover{cursor:pointer}.qwU25c,.qwU25c:hover,.qwU25c:active{color:#7f7f7f;pointer-events:none;opacity:0.5}.FJJygb,.Z3WPhc,.LhKRUe{-moz-box-sizing:border-box;box-sizing:border-box}.FJJygb{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-flow:column nowrap;pointer-events:none;position:fixed;width:100%;z-index:1200}.FJJygb.qwLQJ{padding:0 1.5rem}@media (max-width:30rem){.FJJygb.qwLQJ{padding:0 .5rem}}.FJJygb.A2eYae{-moz-box-align:start;align-items:flex-start;bottom:1.5rem;padding:0 1.5rem}.FJJygb.qwLQJ .LhKRUe{margin-bottom:.5rem}.FJJygb.A2eYae .LhKRUe{margin-top:.5rem}.Z3WPhc{pointer-events:auto}.FJJygb.qwLQJ .Z3WPhc{max-width:47.5rem}.FJJygb.A2eYae .Z3WPhc{max-width:35.5rem}.LhKRUe{letter-spacing:.0142857143em;font-family:Roboto,Arial,sans-serif;font-size:.875rem;font-weight:400;line-height:1.25rem;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);-moz-box-align:center;align-items:center;background-color:rgb(32,33,36);border-radius:.25rem;color:rgb(232,234,237);display:-moz-box;display:flex;fill:rgb(232,234,237);-moz-box-pack:justify;justify-content:space-between;min-height:3rem;min-width:21.5rem;padding:.75rem 1rem}.LhKRUe.JKIkqc{background-color:rgb(179,20,18)}.LhKRUe.JKIkqc,.LhKRUe.JKIkqc .eoooNd{color:#fff}.U51CBd{margin-right:1rem}.eoooNd.eoooNd{height:auto;flex-shrink:0;margin-bottom:0;margin-top:0;white-space:nowrap}.ar1wZ{margin:0 -.375rem 0 .75rem}.dzWTB{display:-webkit-box;overflow:hidden;text-overflow:ellipsis;word-break:break-word;-webkit-line-clamp:2;-webkit-box-orient:vertical}.VfPpkd-r7nwK{color:#fff;color:var(--mdc-theme-surface,#fff)}.VfPpkd-r7nwK{background-color:#6200ee;background-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-gkkIFf,.VfPpkd-WLXbod{min-width:344px}@media (max-width:344px),(max-width:480px){.VfPpkd-gkkIFf,.VfPpkd-WLXbod{min-width:100%}}.VfPpkd-gkkIFf{max-width:720px}.VfPpkd-ORHb{z-index:1;border-bottom-style:solid;-moz-box-sizing:border-box;box-sizing:border-box;display:none;flex-shrink:0;height:0;position:relative;width:100%}@media (max-width:480px){.VfPpkd-ORHb .VfPpkd-WLXbod{left:0;right:0}.VfPpkd-ORHb .VfPpkd-Rj7Y9b{margin-left:16px;margin-right:36px}[dir=rtl] .VfPpkd-ORHb .VfPpkd-Rj7Y9b,.VfPpkd-ORHb .VfPpkd-Rj7Y9b[dir=rtl]{margin-left:36px;margin-right:16px}}@media (max-width:480px){.VfPpkd-ORHb.VfPpkd-ORHb-OWXEXe-N4imRe-eu7FSc .VfPpkd-gkkIFf{flex-wrap:wrap}.VfPpkd-ORHb.VfPpkd-ORHb-OWXEXe-N4imRe-eu7FSc .VfPpkd-r7nwK{margin-bottom:12px}.VfPpkd-ORHb.VfPpkd-ORHb-OWXEXe-N4imRe-eu7FSc .VfPpkd-Rj7Y9b{margin-left:16px;margin-right:8px;padding-bottom:4px}[dir=rtl] .VfPpkd-ORHb.VfPpkd-ORHb-OWXEXe-N4imRe-eu7FSc .VfPpkd-Rj7Y9b,.VfPpkd-ORHb.VfPpkd-ORHb-OWXEXe-N4imRe-eu7FSc .VfPpkd-Rj7Y9b[dir=rtl]{margin-left:8px;margin-right:16px}.VfPpkd-ORHb.VfPpkd-ORHb-OWXEXe-N4imRe-eu7FSc .VfPpkd-rfWUU{margin-left:auto}}.VfPpkd-ORHb-OWXEXe-uGFO6d,.VfPpkd-ORHb-OWXEXe-FNFY6c,.VfPpkd-ORHb-OWXEXe-FnSee{display:-moz-box;display:flex}.VfPpkd-ORHb-OWXEXe-FNFY6c{transition:height .3s ease}.VfPpkd-ORHb-OWXEXe-FNFY6c .VfPpkd-gkkIFf{transition:transform .3s ease;transform:translateY(0)}.VfPpkd-ORHb-OWXEXe-FnSee{transition:height .25s ease}.VfPpkd-ORHb-OWXEXe-FnSee .VfPpkd-gkkIFf{transition:transform .25s ease}.VfPpkd-ORHb-OWXEXe-VErWse .VfPpkd-gkkIFf{left:0;margin-left:auto;margin-right:auto;right:0}.VfPpkd-WLXbod{border-bottom-style:solid;-moz-box-sizing:border-box;box-sizing:border-box;height:inherit;position:fixed;width:100%}.VfPpkd-gkkIFf{display:-moz-box;display:flex;min-height:52px;position:absolute;transform:translateY(-100%);width:100%}.VfPpkd-r7nwK-fmcmS-sM5MNb{display:-moz-box;display:flex;width:100%}.VfPpkd-r7nwK{margin-left:16px;margin-right:0;flex-shrink:0;margin-top:16px;margin-bottom:16px;text-align:center}[dir=rtl] .VfPpkd-r7nwK,.VfPpkd-r7nwK[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-w255rc{position:relative;top:50%;transform:translateY(-50%)}.VfPpkd-Rj7Y9b{margin-left:24px;margin-right:90px;align-self:center;-moz-box-flex:1;flex-grow:1;padding-top:16px;padding-bottom:16px}[dir=rtl] .VfPpkd-Rj7Y9b,.VfPpkd-Rj7Y9b[dir=rtl]{margin-left:90px;margin-right:24px}.VfPpkd-rfWUU{padding-left:0;padding-right:8px;align-self:flex-end;display:-moz-box;display:flex;flex-shrink:0;padding-bottom:8px;padding-top:8px}[dir=rtl] .VfPpkd-rfWUU,.VfPpkd-rfWUU[dir=rtl]{padding-left:8px;padding-right:0}.VfPpkd-ORHb{background-color:#fff;background-color:var(--mdc-banner-container-color,#fff);border-bottom-color:rgba(0,0,0,.12);border-bottom-color:var(--mdc-banner-divider-color,rgba(0,0,0,.12));border-bottom-width:1px;border-bottom-width:var(--mdc-banner-divider-height,1px);border-radius:0;border-radius:var(--mdc-banner-container-shape,0)}.VfPpkd-ORHb .VfPpkd-Rj7Y9b{color:#000;color:var(--mdc-banner-supporting-text-color,#000)}.VfPpkd-ORHb .VfPpkd-Rj7Y9b{letter-spacing:.0178571429em;letter-spacing:var(--mdc-banner-supporting-text-tracking,.0178571429em);font-size:.875rem;font-size:var(--mdc-banner-supporting-text-size,.875rem);font-family:Roboto,sans-serif;font-family:var(--mdc-banner-supporting-text-font,Roboto,sans-serif);font-weight:400;font-weight:var(--mdc-banner-supporting-text-weight,400);line-height:1.25rem;line-height:var(--mdc-banner-supporting-text-line-height,1.25rem)}.VfPpkd-ORHb .VfPpkd-r7nwK{border-radius:50%;border-radius:var(--mdc-banner-with-image-image-shape,50%)}.VfPpkd-ORHb .VfPpkd-r7nwK{height:40px;height:var(--mdc-banner-with-image-image-size,40px);width:40px;width:var(--mdc-banner-with-image-image-size,40px)}.VfPpkd-ORHb .VfPpkd-WLXbod{background-color:#fff;background-color:var(--mdc-banner-container-color,#fff)}.VfPpkd-ORHb .VfPpkd-WLXbod{border-bottom-color:rgba(0,0,0,.12);border-bottom-color:var(--mdc-banner-divider-color,rgba(0,0,0,.12))}.VfPpkd-ORHb .VfPpkd-WLXbod{border-bottom-width:1px;border-bottom-width:var(--mdc-banner-divider-height,1px)}.VfPpkd-ORHb .VfPpkd-LgbsSe:not(:disabled){color:#6200ee;color:var(--mdc-text-button-label-text-color,var(--mdc-banner-action-label-text-color,#6200ee))}.VfPpkd-ORHb .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-ORHb .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{background-color:#6200ee;background-color:var(--mdc-text-button-hover-state-layer-color,var(--mdc-banner-action-hover-state-layer-color,#6200ee))}.VfPpkd-ORHb .VfPpkd-LgbsSe:hover .VfPpkd-Jh9lGc::before,.VfPpkd-ORHb .VfPpkd-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-text-button-hover-state-layer-opacity,var(--mdc-banner-action-hover-state-layer-opacity,.04))}.VfPpkd-ORHb .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-ORHb .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-text-button-focus-state-layer-opacity,var(--mdc-banner-action-focus-state-layer-opacity,.12))}.VfPpkd-ORHb .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-ORHb .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-text-button-pressed-state-layer-opacity,var(--mdc-banner-action-pressed-state-layer-opacity,.1))}.VfPpkd-ORHb .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-text-button-pressed-state-layer-opacity,var(--mdc-banner-action-pressed-state-layer-opacity,0.1))}.VfPpkd-jsLfKf-JIbuQc{margin-left:0;margin-right:8px}[dir=rtl] .VfPpkd-jsLfKf-JIbuQc,.VfPpkd-jsLfKf-JIbuQc[dir=rtl]{margin-left:8px;margin-right:0}.geqPvd{background-color:#fff;border-bottom-color:rgb(218,220,224)}.geqPvd .VfPpkd-WLXbod{background-color:#fff}.geqPvd .VfPpkd-Rj7Y9b{color:rgb(60,64,67)}.geqPvd .VfPpkd-WLXbod{border-bottom-color:rgb(218,220,224)}.geqPvd .VfPpkd-r7nwK{color:#fff}.geqPvd .VfPpkd-r7nwK{background-color:rgb(26,115,232)}.geqPvd .VfPpkd-LgbsSe:not(:disabled){background-color:transparent}.geqPvd .VfPpkd-LgbsSe:not(:disabled){color:rgb(26,115,232);color:var(--gm-colortextbutton-ink-color,rgb(26,115,232))}.geqPvd .VfPpkd-LgbsSe:disabled{color:rgba(60,64,67,.38);color:var(--gm-colortextbutton-disabled-ink-color,rgba(60,64,67,.38))}.geqPvd .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.geqPvd .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.geqPvd .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.geqPvd .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.geqPvd .VfPpkd-LgbsSe:hover:not(:disabled),.geqPvd .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.geqPvd .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.geqPvd .VfPpkd-LgbsSe:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-colortextbutton-ink-color--stateful,rgb(23,78,166))}.geqPvd .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.geqPvd .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-colortextbutton-state-color,rgb(26,115,232))}.geqPvd .VfPpkd-LgbsSe:hover .VfPpkd-Jh9lGc::before,.geqPvd .VfPpkd-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.geqPvd .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.geqPvd .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.geqPvd .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.geqPvd .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.geqPvd .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.geqPvd .UMrnmb-jsLfKf-JIbuQc{margin-right:8px}.skamq{background-color:rgb(179,20,18)}.neGRTd #gb{font-family:"Roboto",Helvetica,Arial,sans-serif;min-width:0!important;padding-right:1.5rem;position:static}@media not all and (max-width:40em){#gbsfw{position:fixed}}.xHPsid{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;justify-content:center;max-width:100%;white-space:nowrap}.xHPsid .hN1OOc{height:4rem}.x1qYbe>.xHPsid{justify-content:normal;padding-left:3.5rem}.TeZa2e{overflow:-moz-scrollbars-none;overflow-x:hidden;overflow-y:hidden}.x1qYbe.TeZa2e{overflow-x:scroll}.QTigq .TeZa2e::-webkit-scrollbar{background:transparent;height:0}.wZTANe{flex-shrink:0;height:100%}.hN1OOc{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;border-bottom:solid 0.125rem transparent;box-sizing:border-box;height:100%;padding:0.125rem 1.5rem 0 1.5rem;position:relative;text-decoration:none}.hN1OOc.eumXzf:after{border-top-width:0.25rem;border-top-style:solid;-moz-border-radius:0.25rem 0.25rem 0 0;border-radius:0.25rem 0.25rem 0 0;bottom:-0.125rem;content:"";height:0;left:0;position:absolute;right:0}@media (max-width:40em){.hN1OOc{padding:0.125rem 1rem 0 1rem}}.hN1OOc:hover,.J1raN:hover{cursor:pointer}.wZTANe .J1raN{color:#5f6368;border-bottom:none;padding-top:0}.wZTANe .J1raN:hover{color:#202124}.mhCMAe{flex-shrink:0;height:4.0625rem}@media (max-width:65.125em){.mwJvDe .ECPFEb{flex-shrink:0;padding-top:4rem}.Xqnlu:not(.QTigq) .ECPFEb{padding-top:5rem}}.Hwv4mb,.Hwv4mb .OGhwGf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;justify-content:center;max-width:100%;overflow:hidden}.Hwv4mb .OGhwGf:focus .Pce5Kb,.Hwv4mb .OGhwGf:hover .Pce5Kb{color:currentcolor}.s7ovNb{padding-top:0.625rem}.joJglb{background:white;border-bottom:0.0625rem solid #e0e0e0;flex-shrink:0;line-height:1.7em;position:fixed;top:0;transform:none;transition:transform cubic-bezier(0.4,0,0.2,1) 240ms;width:100%;z-index:986}.joJglb.yeBmWb{transform:translateY(calc(-100% - 0.5rem*1))}.yeBmWb .FJJygb.qwLQJ{margin-top:0.5rem}.joJglb.kLHn3{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15)}.XIpEib{height:4rem;padding-left:1.5rem}.R2tE8e{justify-content:center;height:4rem;padding-right:1rem;text-align:center;width:100%}.Mtd4hb{justify-content:flex-end;flex-shrink:0;padding-right:0.5rem}.kWv2Xb{flex-shrink:0;height:1.5rem}.XGLVqf{margin-right:1rem}.PYWmSe{flex-shrink:0;margin-right:-moz-calc(-36px + 1rem*1);margin-right:calc(-36px + 1rem*1);margin-left:-moz-calc(-48px + 1rem*1);margin-left:calc(-48px + 1rem*1)}.aTtRxf{bottom:0;position:absolute;left:0;right:0}.k43Owe{flex-shrink:0;margin-right:1rem}.AMagsb:after{color:red;content:"FakeRubricsEnabled";display:block}@media not all and (max-width:65.125em){.meR3Qc{display:none}.FXKA9c,.Mtd4hb{-moz-box-flex:1 1 0.0625rem;flex:1 1 0.0625rem;min-width:0}.R2tE8e{margin:0 1rem;width:auto}}@media (max-width:65.125em){.VHRSDf{display:none}.FXKA9c{box-flex:1;flex-grow:1;min-width:0;overflow:hidden;margin-right:1rem}}.fXYYpf{display:-moz-box;display:flex}.fXYYpf .T4LgNb{display:block;-moz-box-flex:1;flex:1 1 auto;min-width:0;position:relative}.T4LgNb{bottom:0;left:0;top:0;right:0;z-index:1}.QMEh5b{top:0;left:0;right:0;z-index:3}.AOq4tb{height:56px}.kFwPee{position:relative;z-index:1}.ydMMEb{height:56px;width:100%}.SSPGKf{overflow-y:hidden;bottom:0;left:0;right:0;top:0}.ecJEib .AOq4tb,.ecJEib .ydMMEb{height:64px}.e2G3Fb.EWZcud .AOq4tb,.e2G3Fb.EWZcud .ydMMEb{height:48px}.e2G3Fb.b30Rkd .AOq4tb,.e2G3Fb.b30Rkd .ydMMEb{height:56px}.SSPGKf{position:relative;min-height:100%}.SSPGKf.BIIBbc{height:100%;overflow:hidden}.kFwPee{backface-visibility:hidden;min-height:100%;height:auto}.T4LgNb{min-height:100%;position:relative}.T4LgNb.eejsDc{min-height:100%;overflow-y:hidden}.QMEh5b{position:fixed}[dir=rtl] .DnNMBb,[dir=rtl] .o1Sh5{transform:scaleX(-1)}.gMIble{background-image:url(data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIHdpZHRoPSIyMzYiIGhlaWdodD0iNzAiIHByZXNlcnZlQXNwZWN0UmF0aW89Im5vbmUiPjxwYXRoIGZpbGw9Im5vbmUiIGQ9Ik0tNDA2LTE0NjRIOTk0djM2MDBILTQwNnoiLz48cGF0aCBkPSJNMjMxIDV2MTRoLTE0VjVoMTRtMC0yaC0xNGMtMS4xIDAtMiAuOS0yIDJ2MTRjMCAxLjEuOSAyIDIgMmgxNGMxLjEgMCAyLS45IDItMlY1YzAtMS4xLS45LTItMi0yeiIvPjxwYXRoIGZpbGw9Im5vbmUiIGQ9Ik0yMTIgMGgyNHYyNGgtMjR6Ii8+PHBhdGggZmlsbD0ibm9uZSIgZD0iTS00MDYtMTA0MEg5OTR2MzYwMEgtNDA2eiIvPjxwYXRoIGZpbGw9Im5vbmUiIGQ9Ik0yMTIgNDBoMjR2MjRoLTI0eiIvPjxwYXRoIGQ9Ik0yMzEgNDNoLTE0Yy0xLjEgMC0yIC45LTIgMnYxNGMwIDEuMS45IDIgMiAyaDE0YzEuMSAwIDItLjkgMi0yVjQ1YzAtMS4xLS45LTItMi0yem0tOSAxNGwtNS01IDEuNC0xLjQgMy42IDMuNiA3LjYtNy42TDIzMSA0OGwtOSA5eiIvPjxnPjxwYXRoIGZpbGwtb3BhY2l0eT0iLjA5IiBkPSJNMCAwaDEwNXY3MEgweiIvPjxwYXRoIGQ9Ik01Mi41IDE1Yy0xMSAwLTIwIDktMjAgMjBzOSAyMCAyMCAyMCAyMC05IDIwLTIwLTktMjAtMjAtMjB6bS0yIDM1LjljLTcuOS0xLTE0LTcuNy0xNC0xNS45IDAtMS4yLjItMi40LjQtMy42bDkuNiA5LjZ2MmMwIDIuMiAxLjggNCA0IDR2My45em0xMy44LTUuMWMtLjUtMS42LTItMi44LTMuOC0yLjhoLTJ2LTZjMC0xLjEtLjktMi0yLTJoLTEydi00aDRjMS4xIDAgMi0uOSAyLTJ2LTRoNGMyLjIgMCA0LTEuOCA0LTR2LS44YzUuOSAyLjQgMTAgOC4xIDEwIDE0LjggMCA0LjItMS42IDcuOS00LjIgMTAuOHoiIGZpbGw9IiNmZmYiLz48L2c+PGc+PHBhdGggZmlsbC1vcGFjaXR5PSIuMDkiIGQ9Ik0xMDYgMGgxMDV2NzBIMTA2eiIvPjxwYXRoIGQ9Ik0xNzMgMjEuMmMtMS4xLS40LTcuOC0uNy0xNC41LS43cy0xMy40LjQtMTQuNS43Yy0yLjguOS0zLjYgNy4yLTMuNiAxMy44cy44IDEyLjkgMy42IDEzLjhjMS4xLjQgNy44LjcgMTQuNS43czEzLjQtLjQgMTQuNS0uN2MyLjgtLjkgMy42LTcuMiAzLjYtMTMuOHMtLjgtMTIuOS0zLjYtMTMuOHptLTE4LjEgMjJWMjYuOGwxMC45IDguMi0xMC45IDguMnoiIGZpbGw9IiNmZmYiLz48L2c+PGc+PHBhdGggZD0iTTIyMS42MjUgMzEuOTdjMC0xLjA1LS41ODMtMS45MjQtMS40NTgtMi4zMzJ2MS4yODRsMS40NTggMS40NTh2LS40MXptMS40NTggMGMwIC41MjYtLjExNiAxLjA1LS4yOTEgMS41MThsLjg3NS44NzVjLjQwOC0uNy41ODMtMS41NzUuNTgzLTIuNDVhNS4yNTkgNS4yNTkgMCAwMC00LjA4My01LjEzM3YxLjIyNWMxLjY5MS41ODMgMi45MTYgMi4wOTkgMi45MTYgMy45NjZ6bS04LjU3NS01LjI1bC0uNzU4Ljc1OSAyLjc0MiAyLjc0MmgtMi43NDJ2My41aDIuMzMzTDIxOSAzNi42Mzh2LTMuOTA5bDIuNTA4IDIuNTA5YTQuODU5IDQuODU5IDAgMDEtMS4zNDEuN3YxLjIyNWE0Ljk2OSA0Ljk2OSAwIDAwMi4xNTgtMS4wNWwxLjE2NyAxLjE2Ny43NTgtLjc1OS01LjI1LTUuMjUtNC40OTItNC41NXptNC40OTIuNTg0bC0xLjIyNSAxLjIyNUwyMTkgMjkuNzU0di0yLjQ1eiIgZmlsbD0iI2RhNDMzNiIvPjxwYXRoIGZpbGw9Im5vbmUiIGQ9Ik0yMTIgMjVoMTR2MTRoLTE0eiIvPjwvZz48L3N2Zz4=);background-repeat:no-repeat;background-size:14.75rem 4.375rem;flex-shrink:0}.N6Z5Rb{background-position:-13.25rem -2.5rem;height:1.5rem;width:1.5rem}.pu837b{background-position:-13.25rem 0;height:1.5rem;width:1.5rem}.aV1rJe{background-position:0 0;height:4.375rem;width:6.5625rem}.dxO7bc{background-position:-6.625rem 0;height:4.375rem;width:6.5625rem}.DnNMBb{background-position:-13.25rem -1.5625rem;height:0.875rem;width:0.875rem}.a6pJXc{display:none}.mIM26c .a6pJXc{display:block}.SRIM0d .Y5vSD,.SRIM0d .nforOe,.SRIM0d .D0cJPb,.SRIM0d .CG2qQ,.SRIM0d .dRIMEd,.SRIM0d .MyrTyc,.SRIM0d .DJd7Z,.SRIM0d .eDpnVe,.SRIM0d .Iz6rbe,.SRIM0d .GKAvYc,.SRIM0d .Nvl44e,.SRIM0d .CMmBPd,.SRIM0d .faqTte,.SRIM0d .nmFHZb,.CPYzFb .Y5vSD,.hhj3ub .nforOe,.nTrDbc .D0cJPb,.Y0qupd .CG2qQ,.MAdsVd .dRIMEd,.GAP4ve .MyrTyc,.MAdsVd.xSXax .DCIKCc,.GAP4ve .TgX6fb,.OYpLJd .TgX6fb,.JL2pRe .Gh0umc,.TIunU .P354se,.nGmYJe .kpDQ8,.AJlUyd .Iz6rbe,.dLNT1b .GKAvYc,.V7D6ud .Nvl44e,.AEGTVe .CMmBPd,.fKVgu .faqTte,.KiTHSb .nmFHZb,.gyaw1d .zzAqTb,.kU4uPd .r8KdYe,.iJzZke .Jp15We,.iJzZke .J2Cevf,.z7HEHd .Jp15We,.Qqqlwf .J2Cevf,.Hlw1k .mmOZjd,.We03Jb .sEZiv,.W0dUmf .GR7QId,.xzRrDe .XztFzd,.OOnEBd>:not(.sH2L2e):not(.xgkURe),.juWHme .Q6ApZc,.mIM26c .YHNy6b,[aria-expanded="true"] .HbKQLd,[aria-expanded="false"] .sjxkNc{display:none;margin:0}@media (max-width:40em){.pOf0gc{display:none!important}}@media (max-width:30em){.nk6WKe .Oe4zIb{display:none;margin:0}}@media not all and (max-width:40em){.nQaZq{display:none!important}}@media (max-width:30em){.EvT0id{display:none!important}}@media not all and (max-width:30em){.Tckeqf{display:none!important}}.hRUMVb{display:inline-block;position:relative;width:32px;height:32px}.eZj3ab{position:absolute;width:0;height:0;overflow:hidden}.EjqBzf{width:100%;height:100%}.hRUMVb.qs41qe .EjqBzf{animation:spinner-container-rotate 1568ms linear infinite}.xgjrdc{position:absolute;width:100%;height:100%;opacity:0}.W16UYe{border-color:#1a73e8}.Z3wgcd{border-color:#d93025}.YAHIzf{border-color:#f9ab00}.zd0Iye{border-color:#1e8e3e}.hRUMVb.qs41qe .xgjrdc.W16UYe{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-blue-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.hRUMVb.qs41qe .xgjrdc.Z3wgcd{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-red-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.hRUMVb.qs41qe .xgjrdc.YAHIzf{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-yellow-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.hRUMVb.qs41qe .xgjrdc.zd0Iye{animation:spinner-fill-unfill-rotate 5332ms cubic-bezier(0.4,0,0.2,1) infinite both,spinner-green-fade-in-out 5332ms cubic-bezier(0.4,0,0.2,1) infinite both}.lUa73{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;top:0;left:45%;width:10%;height:100%;overflow:hidden;border-color:inherit}.lUa73 .O8fgAf{width:1000%;left:-450%}.NzjLhf{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;top:0;width:50%;height:100%;overflow:hidden;border-color:inherit}.NzjLhf.GBKMJf{left:0}.NzjLhf.W8OIte{left:50%}.NzjLhf .O8fgAf{width:200%}.O8fgAf{position:absolute;top:0;right:0;bottom:0;left:0;-moz-box-sizing:border-box;box-sizing:border-box;height:100%;border-width:3px;border-style:solid;border-color:inherit;border-bottom-color:transparent;-moz-border-radius:50%;border-radius:50%;animation:none}.NzjLhf.GBKMJf .O8fgAf{border-right-color:transparent;transform:rotate(129deg)}.NzjLhf.W8OIte .O8fgAf{left:-100%;border-left-color:transparent;transform:rotate(-129deg)}.hRUMVb.qs41qe .NzjLhf.GBKMJf .O8fgAf{animation:spinner-left-spin 1333ms cubic-bezier(0.4,0,0.2,1) infinite both}.hRUMVb.qs41qe .NzjLhf.W8OIte .O8fgAf{animation:spinner-right-spin 1333ms cubic-bezier(0.4,0,0.2,1) infinite both}.hRUMVb.sf4e6b .EjqBzf{animation:spinner-container-rotate 400ms linear infinite,spinner-fade-out 400ms cubic-bezier(0.4,0,0.2,1)}@keyframes spinner-container-rotate{to{transform:rotate(360deg)}}@keyframes spinner-fill-unfill-rotate{12.5%{transform:rotate(135deg)}25%{transform:rotate(270deg)}37.5%{transform:rotate(405deg)}50%{transform:rotate(540deg)}62.5%{transform:rotate(675deg)}75%{transform:rotate(810deg)}87.5%{transform:rotate(945deg)}to{transform:rotate(1080deg)}}@keyframes spinner-blue-fade-in-out{0%{opacity:.99}25%{opacity:.99}26%{opacity:0}89%{opacity:0}90%{opacity:.99}to{opacity:.99}}@keyframes spinner-red-fade-in-out{0%{opacity:0}15%{opacity:0}25%{opacity:.99}50%{opacity:.99}51%{opacity:0}}@keyframes spinner-yellow-fade-in-out{0%{opacity:0}40%{opacity:0}50%{opacity:.99}75%{opacity:.99}76%{opacity:0}}@keyframes spinner-green-fade-in-out{0%{opacity:0}65%{opacity:0}75%{opacity:.99}90%{opacity:.99}to{opacity:0}}@keyframes spinner-left-spin{0%{transform:rotate(130deg)}50%{transform:rotate(-5deg)}to{transform:rotate(130deg)}}@keyframes spinner-right-spin{0%{transform:rotate(-130deg)}50%{transform:rotate(5deg)}to{transform:rotate(-130deg)}}@keyframes spinner-fade-out{0%{opacity:.99}to{opacity:0}}.jsbB5e{-moz-user-select:none;-moz-user-select:none;display:inline-block;outline:none;width:280px}.jsbB5e.mXfoO{width:100%}.Yalane{min-height:1.5em;position:relative;vertical-align:top}.fWf7qe .Yalane{background-color:#f8f9fa;-moz-border-radius:4px 4px 0 0;border-radius:4px 4px 0 0}.fWf7qe.RDPZE .Yalane{background-color:rgba(248,249,250,.38)}.fWf7qe:not(.RDPZE):hover .Yalane{background-color:#f1f3f4;cursor:pointer}.AkVYk .Yalane{-moz-border-radius:4px;border-radius:4px}.Y6Mzcf{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;position:relative}.AkVYk .Yalane:before{border:1px solid #dadce0;-moz-border-radius:4px;border-radius:4px;bottom:0;content:"";left:0;position:absolute;right:0;top:0;z-index:0}.AkVYk.u3bW4e .Yalane:before{border:2px solid #1a73e8}.AkVYk.IYewr .Yalane:before{border:2px solid #d93025}.AkVYk.IYewr.RDPZE .Yalane:before{border:2px solid rgba(217,48,37,.38)}.hqfVKd{box-flex:1;flex-grow:1;flex-shrink:1;font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;background-color:transparent;border:none;-moz-box-sizing:content-box;box-sizing:content-box;caret-color:#1a73e8;display:block;height:24px;min-height:24px;margin:0;outline:none;overflow-y:visible;overflow-x:hidden;padding:16px;resize:none;white-space:pre-wrap;word-wrap:break-word;z-index:1}.jsbB5e.IYewr .hqfVKd{caret-color:#d93025}.jsbB5e.IYewr.RDPZE .hqfVKd{caret-color:rgba(217,48,37,.38)}.fWf7qe:not(.yaevDc) .hqfVKd{padding:23px 16px 9px 16px}.jsbB5e.KoF8Ce .hqfVKd,.fWf7qe.KoF8Ce:not(.yaevDc) .hqfVKd{padding-bottom:0}.fWf7qe.u3bW4e .Yalane,.fWf7qe.CDELXb .Yalane,.fWf7qe.IhU0Je .Yalane{padding-top:23px}.AkVYk.u3bW4e .Yalane,.AkVYk.CDELXb .Yalane,.AkVYk.IhU0Je .Yalane,.jsbB5e.IbzNie.yaevDc .Yalane,.fWf7qe.u3bW4e.yaevDc .Yalane,.fWf7qe.CDELXb.yaevDc .Yalane{padding-top:16px}.jsbB5e.u3bW4e .hqfVKd,.jsbB5e.CDELXb.yaevDc .hqfVKd,.jsbB5e.IbzNie.yaevDc .hqfVKd,.fWf7qe:not(.yaevDc).u3bW4e .hqfVKd,.AkVYk:not(.yaevDc).u3bW4e .hqfVKd,.fWf7qe:not(.yaevDc).CDELXb .hqfVKd,.AkVYk:not(.yaevDc).CDELXb .hqfVKd,.fWf7qe:not(.yaevDc).IhU0Je .hqfVKd,.AkVYk:not(.yaevDc).IhU0Je .hqfVKd{padding-top:0}.hqfVKd.bhfTYe{text-align:center}.jsbB5e.RDPZE .hqfVKd{color:rgba(60,64,67,.38)}.oQ5Hqe{background-color:#80868b;bottom:0;height:1px;left:0;margin:0;padding:0;position:absolute;width:100%}.aCxcAe{-moz-transform:scaleX(0);transform:scaleX(0);background-color:#1a73e8;bottom:0;height:2px;left:0;margin:0;padding:0;position:absolute;width:100%}.fWf7qe.RDPZE .oQ5Hqe{background-color:rgba(128,134,139,.38)}.AkVYk .oQ5Hqe,.AkVYk .aCxcAe{display:none}.jsbB5e.IYewr>.Yalane>.oQ5Hqe,.jsbB5e.IYewr>.Yalane>.aCxcAe{background-color:#d93025;height:2px}.jsbB5e.IYewr.RDPZE>.Yalane>.oQ5Hqe,.jsbB5e.IYewr.RDPZE>.Yalane>.aCxcAe{background-color:rgba(217,48,37,.38)}.jsbB5e .aCxcAe.Y2Zypf{-moz-animation:agmTextInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:agmTextInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1)}.jsbB5e.u3bW4e>.Yalane>.aCxcAe{-moz-animation:agmTextInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:agmTextInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);-moz-transform:scaleX(1);transform:scaleX(1)}.CYSZae{font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;-moz-transform-origin:bottom left;transform-origin:bottom left;-moz-transition:all .3s cubic-bezier(0.4,0,0.2,1);transition:all .3s cubic-bezier(0.4,0,0.2,1);transition-property:color,top,-webkit-transform;transition-property:color,top,transform;transition-property:color,top,transform,-webkit-transform;color:#5f6368;left:16px;overflow:hidden;pointer-events:none;position:absolute;right:16px;text-overflow:ellipsis;top:16px;white-space:nowrap;z-index:2}.fWf7qe.u3bW4e>.Yalane>.CYSZae,.fWf7qe.CDELXb>.Yalane>.CYSZae,.fWf7qe.IhU0Je>.Yalane>.CYSZae{-moz-transform:scale(.75) translateY(-20px);transform:scale(.75) translateY(-20px)}.AkVYk .CYSZae{background-color:white;padding:2px 4px;left:12px;max-width:-moz-calc(100% - 32px);max-width:calc(100% - 32px);top:14px;right:unset}.AkVYk.u3bW4e>.Yalane>.CYSZae,.AkVYk.CDELXb>.Yalane>.CYSZae,.AkVYk.IhU0Je>.Yalane>.CYSZae{-moz-transform:scale(.75) translateY(-41px);transform:scale(.75) translateY(-41px)}.jsbB5e.u3bW4e .CYSZae{color:#1a73e8}.jsbB5e.RDPZE .CYSZae{color:rgba(60,64,67,.38)}.jsbB5e.IYewr .CYSZae,.jsbB5e.u3bW4e.IYewr .CYSZae{color:#d93025}.jsbB5e.RDPZE.IYewr .Yalane .CYSZae{color:rgba(217,48,37,.38)}.sLGmhc{font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;color:#9aa0a6;left:16px;overflow:hidden;pointer-events:none;position:absolute;right:16px;text-overflow:ellipsis;top:16px;white-space:nowrap;z-index:2}.jsbB5e.RDPZE .sLGmhc{color:rgba(154,160,166,.38)}.fWf7qe:not(.yaevDc) .sLGmhc{top:23px}.jsbB5e.CDELXb>.Yalane>.sLGmhc{display:none}.YQwhRe{font-family:Roboto,Arial,sans-serif;font-size:12px;font-weight:400;letter-spacing:.3px;line-height:16px;height:16px;margin-left:auto;padding-bottom:4px;padding-right:16px;pointer-events:none;text-align:right;white-space:nowrap}.jsbB5e.sT3Fhb{padding-bottom:4px}.yJqEpe,.JmRlzf:not(:empty){font-family:Roboto,Arial,sans-serif;font-size:12px;font-weight:400;letter-spacing:.3px;line-height:16px;flex:1 1 auto;min-height:16px;padding:4px 16px}.jsbB5e.sT3Fhb .K7PyWb{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex}.JmRlzf{pointer-events:none;color:#5f6368}.YQwhRe{color:#5f6368}.jsbB5e.RDPZE .JmRlzf,.jsbB5e.RDPZE .YQwhRe{color:rgba(95,99,104,.38)}.yJqEpe{color:#d93025}.jsbB5e.RDPZE .yJqEpe{color:rgba(217,48,37,.38)}.jsbB5e.k0tWj .JmRlzf,.jsbB5e:not(.k0tWj) .JmRlzf:not(:empty)+.yJqEpe{display:none}.fb0g6{position:relative}.dAR2{background:none;box-shadow:none}.dBlsqc{-moz-box-align:stretch;align-items:stretch;max-width:100%;width:280px}.XXjd3c{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;outline:none;text-align:center}.cOzIj{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1.125rem;letter-spacing:0;font-weight:400;color:rgb(60,64,67);margin:8px 0 0;text-align:center}.UzQuCe{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400;color:rgb(60,64,67);margin-top:8px}.wbPDB{width:100%}.Ajv1wf{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-pack:center;justify-content:center}.a7OWub{flex-shrink:0;line-height:0;padding:0.5rem}.a7OWub:focus{background-color:rgba(153,153,153,.4);-moz-border-radius:50%;border-radius:50%;overflow:hidden;transition:background 150ms}.hVNH5c{box-shadow:0 2px 1px -1px rgba(0,0,0,0.2),0 1px 1px 0 rgba(0,0,0,0.141),0 1px 3px 0 rgba(0,0,0,0.122);-moz-border-radius:4px;border-radius:4px;max-width:280px!important}.hVNH5c.llrsB{max-width:none!important}.hVNH5c .K0NPx{max-width:100%;min-width:0!important;padding:8px 0}.hVNH5c.e5Emjc .FeRvI{padding-left:40px}.FeRvI{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:32px;min-width:112px;overflow:hidden;padding:0}.MEhszc .FeRvI{height:48px}.FeRvI.N2RpBe{background-color:rgba(26,115,232,0.039)}.FeRvI.N2RpBe:hover{background-color:rgba(26,115,232,0.078)}.hVNH5c:not(.MEhszc) .FeRvI.N2RpBe::before{top:0}.FeRvI.N2RpBe.RDPZE{background-color:transparent}.FeRvI .oJeWuf{font-family:Roboto,Arial,sans-serif;font-size:14px;font-weight:400;letter-spacing:.1px;box-sizing:border-box;height:32px;line-height:32px;padding:0 16px;width:100%}.MEhszc .FeRvI .oJeWuf{font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;height:48px;line-height:48px}.FeRvI .jO7h3c{text-overflow:ellipsis;overflow:hidden}.FeRvI .Ce1Y1c{bottom:6px;height:20px;width:20px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;left:16px;opacity:1;top:6px}.MEhszc .FeRvI .Ce1Y1c{bottom:0;height:100%;top:0}.FeRvI .HhLEze{padding:0}.Sa0J5{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;width:100%}.Niache{border-right:0.0625rem solid #e0e0e0}.bHOAdb{flex-shrink:0;position:relative}.nGmYJe .bHOAdb{opacity:0.4}.bHOAdb{height:4.375rem;overflow:hidden;width:6.5625rem}.bHOAdb img,.bHOAdb .mXQw7d{box-sizing:border-box;max-height:100%;max-width:100%}.bHOAdb img.csnH7d{padding:0.375rem}.zyJ7l{background-color:#fafafa}.zyJ7l img{max-height:80%}.F4mChd .bHOAdb{height:3.5rem;width:3.5rem}.JkIgWb{text-decoration:none;outline:none}.QDKOcc{text-overflow:ellipsis;overflow:hidden;white-space:nowrap}.kMUPoc .iv7Rwd{display:none}.DHmSPe{margin-right:-0.5rem}.K013Jb{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;margin-top:0.5rem}.bHOAdb:empty{border:0.0625rem solid #e0e0e0;background:#eee}.MlZb9c.JY4wBc:not(:empty),.MlZb9c.Zat4re:not(:empty){margin-bottom:1rem}.MlZb9c.Zat4re .t2wIBc:not(:first-child) .r0VQac,.MlZb9c.Zat4re .Yzgtqe.WKpRFb:not(:first-child){margin-top:0.75rem}.JY4wBc .t2wIBc:not(:first-child) .r0VQac{margin-top:0.5rem}.r0VQac,.Yzgtqe,.M4LFnf{padding-right:0.5rem}.r0VQac{position:relative}.Yzgtqe{position:relative;overflow:visible}.Yzgtqe .bHOAdb{overflow:hidden;-moz-border-radius:0.4375rem 0 0 0.4375rem;border-radius:0.4375rem 0 0 0.4375rem}.r0VQac .lwlIqf,.Yzgtqe .lwlIqf{bottom:0;left:0;position:absolute;right:0}@media not all and (max-width:40em){.luto0c{position:relative}.luto0c .lwlIqf{bottom:0;left:0;position:absolute;right:0}}.r0VQac .F1bQqd,.r0VQac .vwNuXe,.Yzgtqe .F1bQqd,.Yzgtqe .vwNuXe,.luto0c .F1bQqd,.luto0c .vwNuXe{box-flex:1;flex-grow:1;overflow:hidden}.r0VQac .bHOAdb,.Yzgtqe .bHOAdb,.luto0c .bHOAdb,.ZgfM9>*{margin-right:1rem}.r0VQac.F4mChd .bHOAdb,.F4mChd .ZgfM9>*{margin-right:0.5rem}.MM30Lb{overflow:hidden}.WInaFd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.ZgfM9{padding-left:1rem}.F4mChd .ZgfM9{padding-left:0.5rem}.ZgfM9 .mUbCce,.ZgfM9 .Y5FYJe{margin-left:-0.5rem;margin-right:-0.25rem}.gCEqcd{margin-right:0.25rem}.tAQe1b{color:#5f6368}.Yzgtqe.WKpRFb .ZgfM9{flex-shrink:0}@media not all and (max-width:60rem){.TTxyDb{display:none}}@media (max-width:60rem){.rEszjc{display:none}.Yzgtqe.WKpRFb{display:block;padding:1rem;padding-bottom:0.5rem}.Yzgtqe.WKpRFb .F1bQqd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-bottom:0.5rem;overflow:visible}.Yzgtqe.WKpRFb .ZgfM9{display:block;padding:0}.Yzgtqe.WKpRFb .ZgfM9>*{margin-right:0;margin-bottom:0.5rem}.Yzgtqe.WKpRFb .mUbCce{margin-left:0.5rem;margin-right:-0.5rem}}.J9GwTe{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.J9GwTe img,.J9GwTe .DPvwYc{color:rgba(0,0,0,.549);-moz-box-flex:0 0 auto;flex:0 0 auto;font-size:1rem;height:1rem;margin:0.5rem;width:1rem}.J9GwTe .QDKOcc{font-weight:400}.qYQ2Fb:not(:empty){margin-right:-0.5rem}.AgzMgb.qYQ2Fb:not(:empty),.AgzMgb .qYQ2Fb:last-child{margin-bottom:-0.5rem}@media (max-width:40em){.d3aYgd:not(:empty){margin-right:-0.5rem}.AgzMgb.d3aYgd:not(:empty),.AgzMgb .d3aYgd:last-child{margin-bottom:-0.5rem}}.qYQ2Fb,.MlZb9c.xLFtvb,.d3aYgd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;-moz-flex-wrap:wrap;flex-wrap:wrap}.Q1Ykn{margin-bottom:0.5rem;margin-right:0.5rem}@media (max-width:40em){.luto0c{margin-bottom:0.5rem;margin-right:0.5rem}}.MlZb9c.xLFtvb .t2wIBc{box-sizing:border-box;margin-bottom:0.75rem;margin-right:0.75rem;width:calc(50% - 0.75rem)}@media not all and (max-width:30em){.MlZb9c.xLFtvb:not(:empty){margin-right:-0.75rem}.AgzMgb.MlZb9c.xLFtvb:not(:empty),.AgzMgb .MlZb9c.xLFtvb:last-child{margin-bottom:-0.75rem}}@media not all and (max-width:40em){.d3aYgd:not(:empty){margin-right:-0.75rem}.AgzMgb.d3aYgd:not(:empty),.AgzMgb .d3aYgd:last-child{margin-bottom:-0.75rem}.d3aYgd .luto0c{box-sizing:border-box;margin-bottom:0.75rem;margin-right:0.75rem;width:calc(50% - 0.75rem)}}@media (max-width:30em){.MlZb9c.xLFtvb{flex-direction:column;-moz-flex-wrap:nowrap;flex-wrap:nowrap}.MlZb9c.xLFtvb .t2wIBc,.MlZb9c.xLFtvb .r0VQac{box-sizing:border-box;margin-right:0;width:100%}}.VkhHKd{align-items:center;border:0.0625rem solid #e0e0e0;-moz-border-radius:1rem;border-radius:1rem;box-sizing:border-box;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;height:2rem;max-width:14.25rem;overflow:hidden;padding:0.25rem 0.75rem;position:relative;z-index:0}.VkhHKd:hover .DAnlhb{opacity:.08}.VkhHKd:focus .DAnlhb{opacity:.24}.VkhHKd:active .gM4mlb{animation:hrRippleTransform .2s cubic-bezier(0,0,0.2,1) forwards;opacity:.08}.VkhHKd.e7EEH,.VkhHKd.e7EEH:active,.VkhHKd.e7EEH:visited{color:inherit;text-decoration:none}.DAnlhb{background-color:#5f6368;bottom:0;left:0;opacity:0;overflow:hidden;position:absolute;right:0;top:0;z-index:-1}.rzTfPe{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:0 0 auto;flex:0 0 auto;font-size:1.125rem;height:1.125rem;margin-right:0.5rem;justify-content:center;width:1.125rem}.rzTfPe .DPvwYc{font-size:1.125rem}.rzTfPe img{height:1.125rem;width:1.125rem}.F8dn3e{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.VfPpkd-NLUYnc-V67aGc{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);position:absolute;left:0;transform-origin:left top;line-height:1.15rem;text-align:left;text-overflow:ellipsis;white-space:nowrap;cursor:text;overflow:hidden;will-change:transform;transition:transform .15s cubic-bezier(.4,0,.2,1),color .15s cubic-bezier(.4,0,.2,1)}[dir=rtl] .VfPpkd-NLUYnc-V67aGc,.VfPpkd-NLUYnc-V67aGc[dir=rtl]{right:0;left:auto;transform-origin:right top;text-align:right}.VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{cursor:auto}.VfPpkd-NLUYnc-V67aGc-OWXEXe-ztc6md:not(.VfPpkd-NLUYnc-V67aGc-OWXEXe-ZYIfFd-ztc6md-vXpfLb)::after{margin-left:1px;margin-right:0;content:"*"}[dir=rtl] .VfPpkd-NLUYnc-V67aGc-OWXEXe-ztc6md:not(.VfPpkd-NLUYnc-V67aGc-OWXEXe-ZYIfFd-ztc6md-vXpfLb)::after,.VfPpkd-NLUYnc-V67aGc-OWXEXe-ztc6md:not(.VfPpkd-NLUYnc-V67aGc-OWXEXe-ZYIfFd-ztc6md-vXpfLb)[dir=rtl]::after{margin-left:0;margin-right:1px}.VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-106%) scale(.75)}.VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-standard .25s 1}@keyframes mdc-floating-label-shake-float-above-standard{0%{transform:translateX(0) translateY(-106%) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(4%) translateY(-106%) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(-4%) translateY(-106%) scale(.75)}100%{transform:translateX(0) translateY(-106%) scale(.75)}}.VfPpkd-RWgCYc-ksKsZd::before,.VfPpkd-RWgCYc-ksKsZd::after{position:absolute;bottom:0;left:0;width:100%;border-bottom-style:solid;content:""}.VfPpkd-RWgCYc-ksKsZd::before{z-index:1}.VfPpkd-RWgCYc-ksKsZd::after{transform:scaleX(0);opacity:0;z-index:2}.VfPpkd-RWgCYc-ksKsZd-OWXEXe-auswjd::after{transform:scaleX(1);opacity:1}.VfPpkd-RWgCYc-ksKsZd-OWXEXe-JD038d::after{opacity:0}.VfPpkd-RWgCYc-ksKsZd::before{border-bottom-width:1px}.VfPpkd-RWgCYc-ksKsZd::after{border-bottom-width:2px}.VfPpkd-RWgCYc-ksKsZd::after{transition:transform .18s cubic-bezier(.4,0,.2,1),opacity .18s cubic-bezier(.4,0,.2,1)}.VfPpkd-NSFCdd-i5vt6e{display:-moz-box;display:flex;position:absolute;top:0;right:0;left:0;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;max-width:100%;height:100%;text-align:left;pointer-events:none}[dir=rtl] .VfPpkd-NSFCdd-i5vt6e,.VfPpkd-NSFCdd-i5vt6e[dir=rtl]{text-align:right}.VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-NSFCdd-MpmGFe{-moz-box-sizing:border-box;box-sizing:border-box;height:100%;pointer-events:none}.VfPpkd-NSFCdd-MpmGFe{-moz-box-flex:1;flex-grow:1}.VfPpkd-NSFCdd-Ra9xwd{-moz-box-flex:0;flex:0 0 auto;width:auto}.VfPpkd-NSFCdd-i5vt6e .VfPpkd-NLUYnc-V67aGc{display:inline-block;position:relative;max-width:100%}.VfPpkd-NSFCdd-i5vt6e .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{text-overflow:clip}.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:133.3333333333%}.VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd{padding-left:0;padding-right:8px;border-top:none}[dir=rtl] .VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd[dir=rtl]{padding-left:8px;padding-right:0}.VfPpkd-NSFCdd-i5vt6e-OWXEXe-di8rgd-V67aGc .VfPpkd-NSFCdd-Ra9xwd{display:none}.VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-NSFCdd-MpmGFe{border-top:1px solid;border-bottom:1px solid}.VfPpkd-NSFCdd-Brv4Fb{border-left:1px solid;border-right:none;width:12px}[dir=rtl] .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-NSFCdd-Brv4Fb[dir=rtl]{border-left:none;border-right:1px solid}.VfPpkd-NSFCdd-MpmGFe{border-left:none;border-right:1px solid}[dir=rtl] .VfPpkd-NSFCdd-MpmGFe,.VfPpkd-NSFCdd-MpmGFe[dir=rtl]{border-left:1px solid;border-right:none}.VfPpkd-NSFCdd-Ra9xwd{max-width:calc(100% - 24px)}.WagS8{align-items:center;background-color:#f8f9fa;border-bottom:0.0625rem solid #dadce0;padding:0 1rem 0 1.5rem}@media not all and (max-width:30em){.WagS8{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}}.MJkJGd{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-shrink:0;justify-content:flex-end}.DZz2Tb{box-flex:1;flex-grow:1;padding:1rem 0.3125rem 0 0}@media not all and (max-width:30em){.DZz2Tb{padding:1rem 0.3125rem 1rem 0}}.NGTSFf,.yIdZrf{flex-shrink:0;margin-left:0.3125rem}.kKn9Nc{visibility:hidden}.rZXyy.YwNp1:not(.xp2dJ),.rZXyy:not(.u0dx8e):not(.ILo0B):not(.xp2dJ){cursor:pointer}.rZXyy.xp2dJ{cursor:-moz-grabbing;cursor:-webkit-grabbing;cursor:grabbing}li.xp2dJ{list-style:none}.xp2dJ{box-shadow:0 4px 4px 0 rgba(60,64,67,.3),0 8px 12px 6px rgba(60,64,67,.15);z-index:9998}.rZXyy.YwNp1,.rZXyy:not(.u0dx8e):not(.ILo0B):not(.xp2dJ):hover,.rZXyy:not(.u0dx8e):not(.ILo0B):not(.xp2dJ):focus{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15)}.UQ5E0{box-shadow:0 3px 5px -1px rgba(0,0,0,.2),0 6px 10px 0 rgba(0,0,0,.14),0 1px 18px 0 rgba(0,0,0,.12)}.q6oraf{box-shadow:0 3px 5px -1px rgba(0,0,0,.2),0 6px 10px 0 rgba(0,0,0,.14),0 1px 18px 0 rgba(0,0,0,.12)}.q6oraf .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:#000;color:var(--mdc-theme-on-surface,#000)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(95,99,104)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(60,64,67)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#000;color:var(--mdc-theme-on-surface,#000)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#000;color:var(--mdc-theme-on-surface,#000)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}.Kb1iQ{margin:-1rem 0}.Kb1iQ .mUbCce{vertical-align:middle}@media (max-width:48.75rem){.bA8Agd{display:none}}@media (max-width:40rem){.Kb1iQ{display:-moz-box;display:flex;flex-wrap:wrap;-moz-box-pack:end;justify-content:flex-end}}.JryN0e{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-pack:justify;justify-content:space-between}@media not all and (max-width:30rem){.JryN0e{margin-bottom:1rem;margin-top:-.5rem}}.JryN0e .gQGHgb{margin:0}.m6GIOd{margin:0 .5rem;vertical-align:middle}.SRX5Hd{height:48px}.uynmgb{margin:0 1rem;vertical-align:middle}.bzD7fd{margin-top:.5rem;z-index:987}.GjZJab.GjZJab{box-shadow:0 1px 2px 0 rgba(32,33,36,.3),0 2px 6px 2px rgba(32,33,36,.15);height:3rem;margin:0;padding:0 1.25rem 0 1rem;border-radius:99px}.GjZJab.GjZJab .VfPpkd-Jh9lGc{border-radius:99px}@keyframes hrExpandableRowListItemSpacingExpanding{0%{margin-top:0}to{margin-top:1rem}}@keyframes hrExpandableRowListItemContentExpandingNew{0%{height:0;opacity:0}50%{opacity:1}}@keyframes hrExpandableRowListItemSpacingCollapsing{0%{margin-top:1rem}to{margin-top:0}}@keyframes hrExpandableRowListItemContentCollapsing{0%{opacity:1}to{height:0;opacity:0}}.OlXwxf,.u73Apc{box-sizing:border-box}.OlXwxf:not(.xp2dJ) .u73Apc{cursor:pointer}.OlXwxf+.lXuxY,.lXuxY+.OlXwxf{border-top:none;margin-top:1rem}.lXuxY{position:relative}.lXuxY .u73Apc{border-color:#e0e0e0}.lXuxY,.pO6AMc,.PqkECe{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);border-radius:0.5rem;overflow:hidden;border-top:none}.lXuxY .u73Apc,.pO6AMc .u73Apc,.PqkECe .u73Apc{-moz-border-radius:0;border-radius:0}.OlXwxf+.lXuxY .u73Apc,.lXuxY+.OlXwxf .u73Apc{box-sizing:border-box;height:3.8125rem;padding-top:0.0625rem}.u73Apc{align-items:center;border-bottom:0.0625rem solid #e0e0e0;border-color:transparent;box-sizing:border-box;height:3.75rem;position:relative;z-index:0}.OlXwxf .SFCE1b{bottom:0;left:0;position:absolute;right:0;top:0;z-index:-1}.OlXwxf.OlXwxf:not(:first-child):hover .u73Apc,.OlXwxf:hover+.OlXwxf .u73Apc,.OlXwxf:not(:first-child).kKn9Nc .u73Apc,.OlXwxf.kKn9Nc+.OlXwxf .u73Apc{box-sizing:border-box;height:3.8125rem;padding-top:0.0625rem}.OlXwxf.OlXwxf:hover,.OlXwxf:hover+.OlXwxf{border-top:none}.UW3s6d{flex-shrink:1;padding:1rem 1.5rem}.OlXwxf .UW3s6d{max-height:40vh;overflow:auto}.mCb5vb .UW3s6d{max-height:-moz-calc(80vh - 7.5rem);max-height:calc(80vh - 7.5rem);overflow:auto}.mCb5vb{box-sizing:border-box;width:100%;max-width:100%}.mCb5vb .Shk6y{margin:0}.mCb5vb .UYUfn{padding:0}.mCb5vb .df5yGe{padding:0;border-bottom:0.0625rem solid #e0e0e0;position:relative}.VZMpte{box-sizing:border-box;height:3.75rem}.OlXwxf:hover+.OlXwxf:not(.lXuxY):focus-within .u73Apc{z-index:-1}.OlXwxf:not(:first-child).pO6AMc,.pO6AMc+.OlXwxf{animation:hrExpandableRowListItemSpacingExpanding 150ms cubic-bezier(0.4,0,0.2,1);animation-fill-mode:forwards}.OlXwxf:not(:first-child).VoEgAc,.VoEgAc+.OlXwxf{animation:hrExpandableRowListItemSpacingCollapsing 150ms cubic-bezier(0.4,0,0.2,1);animation-fill-mode:forwards}.OlXwxf.VoEgAc+.OlXwxf.pO6AMc,.OlXwxf.VoEgAc+.OlXwxf.lXuxY,.OlXwxf.PqkECe+.OlXwxf.VoEgAc,.OlXwxf.lXuxY+.OlXwxf.VoEgAc,.OlXwxf.pO6AMc+.OlXwxf.VoEgAc{animation:none}.OlXwxf.AZd1I+.OlXwxf.lXuxY{animation:none;transition:margin-top .3s cubic-bezier(0.4,0,0.2,1)}.S9CVKb{box-sizing:border-box}.OlXwxf.pO6AMc .S9CVKb{animation:hrExpandableRowListItemContentExpandingNew 500ms cubic-bezier(0.4,0,0.2,1);overflow:hidden}.OlXwxf.lXuxY .S9CVKb{transition:height .3s cubic-bezier(0.4,0,0.2,1)}.OlXwxf.VoEgAc .S9CVKb{animation:hrExpandableRowListItemContentCollapsing 500ms cubic-bezier(0.4,0,0.2,1);animation-fill-mode:forwards}.VoEgAc .S9CVKb{overflow:hidden}.AZd1I:not(.VoEgAc) .S9CVKb,.zvbGS .S9CVKb{display:none;height:0!important;visibility:hidden}.OlXwxf.PqkECe .S9CVKb{height:0!important;overflow:hidden}.fPotmc,.NCzUzb{padding:0.375rem 0.5rem}.NCzUzb.dDKhVc{color:#d50000}.akrp3c{display:block}.akrp3c .snByac{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:0.75rem;font-weight:400;line-height:1rem;padding-bottom:0.375rem;padding-top:0.375rem}.L4Hgye{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.L4Hgye:not(:empty),.UbHeTc{margin-bottom:-0.25rem}.UbHeTc .e0pgvc{margin-right:0.25rem;padding-bottom:3px;vertical-align:middle}.kRYv9b{margin-right:0.25rem}@media not all and (max-width:60rem){.ii9Rh{display:none}}.sVNOQ{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.KiTkLc{flex-shrink:0}.k3J5ed{flex-shrink:0;font-weight:400;margin-right:0.25rem}.k3J5ed:not(:empty){margin-left:1rem}.k3J5ed>:not(:last-child),.KiTkLc>:not(:last-child){margin-right:0.5rem}.jrOV5e{color:rgba(0,0,0,.42);fill:rgba(0,0,0,.42);font-size:1.25rem}.DodiNb{margin-right:0.25rem}.seqYL{color:rgba(0,0,0,.38);flex-shrink:0;font-size:.75rem;font-weight:500;line-height:.9375rem;margin-left:.5rem}.seqYL .GHykUb{margin-right:.25rem}.VVwgJb{display:-moz-box;display:flex}.qk5dFc{opacity:.001}.wJ76ge .qk5dFc:focus,.wJ76ge:hover .qk5dFc{opacity:1}.pMq3Db{margin-bottom:1rem}.wJ76ge.nGmYJe{opacity:.57}.WqfsMd{height:2rem;margin:.4rem 1rem 0 0;width:2rem}.G0rp{-moz-box-flex:1;flex-grow:1;min-width:0}.YU7iib{display:-moz-box;display:flex;-moz-box-pack:justify;justify-content:space-between;min-height:1.5rem}.gJItbc{display:inline;margin-right:.5rem}.thiSD{display:-moz-box;display:flex;margin-left:.5rem}.VSWCL{word-wrap:break-word}.KYmC8d,.L8jEMd{margin-left:.5rem}.wJ76ge .a7OWub{padding:0}.q9pD9{border-bottom:.0625rem solid rgb(218,220,224);border-top:.0625rem solid rgb(218,220,224);margin-bottom:1rem;padding:1rem 0 .5rem}.BQa3Cf{-moz-box-flex:1;flex-grow:1}.iS4pCd{margin:1rem 0}.pYglbf .uArJ5e:not(:last-child){margin-right:1rem}.pYglbf .EmVfjc{height:1.125rem;margin:.05625rem;width:1.125rem}@media (max-width:40rem){.XAoEbc .BQa3Cf{margin-top:0}}.PeGHgb.jbH5ac{margin:-1rem -1.5rem}.PeGHgb.Q8U8uc .amzDAb,.PeGHgb:not(.Q8U8uc) .WuChGe,.PeGHgb:not(.Q8U8uc) .VYv8If{display:none}.yoORU{border-bottom:0.0625rem solid #e0e0e0;flex-direction:column;box-flex:1;flex-grow:1;padding:1.5rem}.FfZdze{align-self:flex-start;margin-bottom:1rem}.fKCeB{background:url('https://www.gstatic.com/classroom/empty_states_comments.png') center no-repeat;background-size:contain;flex-shrink:0;height:9rem;margin-bottom:1.5rem;width:9rem}.PeGHgb .f0kHoc{margin:1.5rem;width:initial}.WuChGe{padding:1rem 1.5rem}.VYv8If{padding:1rem 0.25rem}.Ono85c{padding:0 1.5rem}.ruTJle{padding:0}.oh9CFb{padding:0 0.5rem 1rem 1.5rem}.fETHd{padding:0 0.5rem 1rem 0}.QGMq0d{padding:1rem 1.5rem}.XNP4U{padding:1rem 1.5rem 1rem 0}.ho6Zoe{margin-right:0.5rem}.xAiME{box-sizing:border-box;display:inline-block;-moz-flex-wrap:wrap;flex-wrap:wrap;line-height:1.5rem;margin-top:0.25rem;padding:0.5rem 0;word-wrap:break-word}.PeGHgb:not(.Q8U8uc) .Ono85c+.oh9CFb,.PeGHgb:not(.Q8U8uc) .ruTJle+.fETHd{padding-top:1rem}.PeGHgb.Q8U8uc .Ono85c+.QGMq0d,.PeGHgb.Q8U8uc .ruTJle+.XNP4U{border-top:0.0625rem solid #e0e0e0}.PeGHgb.jbH5ac .QGMq0d,.PeGHgb.jbH5ac .XNP4U{margin-left:1.5rem;margin-right:1.5rem;padding-left:0;padding-right:0}.PeGHgb[aria-expanded="false"] .dZVZab:not(:last-child){display:none}.PeGHgb.YHeUvc[aria-expanded="false"] .Ono85c,.PeGHgb.YHeUvc.Q8U8uc[aria-expanded="false"] .oh9CFb,.PeGHgb.YHeUvc.Q8U8uc[aria-expanded="false"] .fETHd,.PeGHgb.YHeUvc.Q8U8uc[aria-expanded="false"] .QGMq0d,.PeGHgb.YHeUvc.Q8U8uc[aria-expanded="false"] .XNP4U{display:none}.A4OZlf{max-width:47.5rem;width:100%}.A4OZlf .wnIM7{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;margin-top:-8px;overflow:auto;padding:8px 0 0 0}.LhPqk .oxacD{display:inline-block}.HM4nYe{width:100%}.isPo5c{display:inline;width:100%}.zJKIV{-moz-user-select:none;-moz-transition:border-color .2s cubic-bezier(0.4,0,0.2,1);transition:border-color .2s cubic-bezier(0.4,0,0.2,1);-moz-border-radius:3px;border-radius:3px;-moz-box-sizing:content-box;box-sizing:content-box;cursor:pointer;display:inline-block;height:20px;outline:none;position:relative;vertical-align:middle;width:20px;z-index:0}.SCWude{-moz-animation:quantumWizPaperAnimateSelectOut .2s forwards;animation:quantumWizPaperAnimateSelectOut .2s forwards;position:relative;width:20px;height:20px;cursor:pointer}[aria-checked=true]>.SCWude{-moz-animation:quantumWizPaperAnimateSelectIn .2s .1s forwards;animation:quantumWizPaperAnimateSelectIn .2s .1s forwards}.t5nRo{position:absolute;top:0;left:0;width:16px;height:16px;-moz-border-radius:50%;border-radius:50%;border:solid 2px;border-color:rgba(0,0,0,.54)}.N2RpBe .t5nRo{border-color:#009688}.wEIpqb{position:absolute;top:50%;left:50%;-moz-border-radius:50%;border-radius:50%;border:5px solid #009688;transition:-webkit-transform ease .28s;transition:transform ease .28s;transition:transform ease .28s,-webkit-transform ease .28s;transform:translateX(-50%) translateY(-50%) scale(0)}[aria-checked=true] .wEIpqb{transform:translateX(-50%) translateY(-50%) scale(1)}.zJKIV[aria-disabled=true]{cursor:default;pointer-events:none}[aria-disabled=true][aria-checked=true] .wEIpqb{border-color:rgba(0,0,0,.26)}[aria-disabled=true] .t5nRo{border-color:rgba(0,0,0,.26)}.k5cvGe{-moz-transform:scale(3);transform:scale(3);-moz-transition:opacity 0.15s ease;transition:opacity 0.15s ease;background-color:rgba(0,0,0,0.2);-moz-border-radius:100%;border-radius:100%;height:20px;left:0;opacity:0;outline:.1px solid transparent;pointer-events:none;position:absolute;width:20px;z-index:-1}.qs41qe>.k5cvGe{-moz-animation:quantumWizRadialInkSpread .3s;animation:quantumWizRadialInkSpread .3s;animation-fill-mode:forwards;opacity:1}.i9xfbb>.k5cvGe{background-color:rgba(0,150,136,0.2)}.u3bW4e>.k5cvGe{-moz-animation:quantumWizRadialInkFocusPulse .7s infinite alternate;animation:quantumWizRadialInkFocusPulse .7s infinite alternate;background-color:rgba(0,150,136,0.2);opacity:1}@keyframes quantumWizPaperAnimateSelectIn{0%{height:0;width:0}to{height:100%;width:100%}}@keyframes quantumWizPaperAnimateSelectOut{0%{height:0;width:0}to{height:100%;width:100%}}.lLfZXe{padding:8px 0}.H2Gmcc{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;align-items:flex-start;flex-direction:column}.lLfZXe.hpDt6e .H2Gmcc{flex-direction:row}.d7L4fc{display:inline-block;flex-shrink:0;height:20px;position:relative;vertical-align:middle;width:20px;z-index:0}.Od2TWd{bottom:-10px;left:-10px;position:absolute;right:-10px;top:-10px;-moz-transition:border-color .2s cubic-bezier(0.4,0,0.2,1);transition:border-color .2s cubic-bezier(0.4,0,0.2,1);-moz-user-select:none;-moz-border-radius:3px;border-radius:3px;box-sizing:border-box;cursor:pointer;height:40px;outline:none;width:40px;z-index:0}.Od2TWd:not(.RDPZE):hover .x0k1lc,.NtlN8c:hover .Od2TWd:not(.RDPZE) .x0k1lc{-moz-transform:scale(2);transform:scale(2);background-color:rgba(26,115,232,0.039);opacity:1}.lLfZXe:not(.hpDt6e) .d7L4fc+.d7L4fc,.lLfZXe:not(.hpDt6e) .NtlN8c+.NtlN8c{margin-top:8px}.lLfZXe.hpDt6e .d7L4fc+.d7L4fc,.lLfZXe.hpDt6e .NtlN8c+.NtlN8c{margin-left:16px}.lLfZXe:not(.x6g5Cd) .d7L4fc+.hHhDYc{margin-left:14px}.NtlN8c{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;align-items:center}.lLfZXe.x6g5Cd .NtlN8c{flex-direction:column-reverse}.hHhDYc{font-family:Roboto,Arial,sans-serif;font-size:16px;font-weight:400;letter-spacing:.1px;line-height:24px;word-break:break-word}.lLfZXe.x6g5Cd .hHhDYc{margin-bottom:8px}.vd3tt{-moz-animation:agmAnimateSelectOut .2s forwards;animation:agmAnimateSelectOut .2s forwards;cursor:pointer;height:20px;position:relative;width:20px}.Od2TWd.N2RpBe>.vd3tt{-moz-animation:agmAnimateSelectIn .2s .1s forwards;animation:agmAnimateSelectIn .2s .1s forwards}.AB7Lab{bottom:10px;left:10px;position:absolute;right:10px;top:10px;border:solid 2px;border-color:#5f6368;-moz-border-radius:50%;border-radius:50%;box-sizing:border-box;height:20px;width:20px}.Od2TWd.N2RpBe .AB7Lab{border-color:#1a73e8}.rseUEf{border:5px solid #1a73e8;-moz-border-radius:50%;border-radius:50%;left:50%;position:absolute;top:50%;transition:-webkit-transform ease .28s;transition:transform ease .28s;transform:translateX(-50%) translateY(-50%) scale(0)}.Od2TWd.N2RpBe .rseUEf{transform:translateX(-50%) translateY(-50%) scale(1)}.Od2TWd.RDPZE{cursor:default;pointer-events:none}.Od2TWd.RDPZE.N2RpBe .rseUEf,.Od2TWd.RDPZE .AB7Lab{border-color:#bdc1c6}.x0k1lc{bottom:10px;left:10px;position:absolute;right:10px;top:10px;-moz-transform:scale(1);transform:scale(1);-moz-transition:opacity .15s ease;transition:opacity .15s ease;background-color:rgba(218,220,224,0.2);-moz-border-radius:100%;border-radius:100%;height:20px;opacity:0;outline:.1px solid transparent;pointer-events:none;width:20px;z-index:-1}.Od2TWd.qs41qe>.x0k1lc{-moz-animation:agmRadialInkSpread .3s;animation:agmRadialInkSpread .3s;animation-fill-mode:forwards;opacity:1}.Od2TWd.u3bW4e>.x0k1lc{-moz-transform:scale(2);transform:scale(2);background-color:rgba(26,115,232,0.122);opacity:1}@keyframes agmRadialInkSpread{0%{-moz-transform:scale(1);transform:scale(1);opacity:0}to{-moz-transform:scale(2);transform:scale(2);opacity:1}}@keyframes agmAnimateSelectIn{0%{height:0;width:0}to{height:100%;width:100%}}@keyframes agmAnimateSelectOut{0%{height:0;width:0}to{height:100%;width:100%}}.rWPWSc{width:20px}.egSPhb .zJKIV,.egSPhb .aMXfFd.bJNwt,.rWPWSc{flex-shrink:0;margin-bottom:0.5rem;margin-right:1rem}.tdmcrb .zJKIV,.tdmcrb .aMXfFd.bJNwt{flex-shrink:0;margin-right:1rem}.JdGGFd,.lbWVCe{background-color:#f1f3f4}.gObdT{box-flex:1;flex-grow:1;justify-content:space-between;margin-bottom:0.5rem;padding:0.5rem 1rem;position:relative;white-space:pre-wrap}.NKFbCb{-moz-border-radius:0.25rem;border-radius:0.25rem}.gObdT.z7tTkd{font-weight:500}.gObdT div{z-index:2}.gObdT .hrBMf{height:100%;left:0;top:0;width:100%;z-index:1}.gObdT .h0pqq{height:100%;left:0;position:absolute;top:0;z-index:0}.LdMiEd .h0pqq{opacity:.08}.lbWVCe .h0pqq{background-color:#dadce0}.EijSib{transition:box-shadow 280ms cubic-bezier(0.4,0,0.2,1);-moz-user-select:none;border:0;-moz-border-radius:16px;border-radius:16px;display:inline-block;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:14px;font-weight:500;letter-spacing:.25px;line-height:36px;text-decoration:none;text-transform:none;line-height:18px;min-width:auto;outline:none;overflow:hidden;position:relative;text-align:center;transition:background .2s .1s;z-index:0}.EijSib:not(.RDPZE){cursor:pointer}.EijSib.qs41qe{transition:box-shadow 280ms cubic-bezier(0.4,0,0.2,1)}.EijSib.RDPZE{color:rgba(0,0,0,.38);fill:rgba(0,0,0,.38)}.kzYc3e.RDPZE{color:rgba(255,255,255,.38);fill:rgba(255,255,255,.38)}.RpYYWb{background-color:#fff;border:1px #dadce0 solid;box-sizing:border-box;color:#3c4043;fill:#3c4043;height:32px}.RpYYWb.qs41qe{box-shadow:0 2px 1px -1px rgba(60,64,67,0.2),0 1px 1px 0 rgba(60,64,67,0.141),0 1px 3px 0 rgba(60,64,67,0.122);border:none;padding:1px}.kzYc3e{background-color:#202124;border:1px #5f6368 solid;color:#f1f3f4;fill:#f1f3f4}.kzYc3e.qs41qe{box-shadow:0 2px 1px -1px rgba(0,0,0,0.2),0 1px 1px 0 rgba(0,0,0,0.141),0 1px 3px 0 rgba(0,0,0,0.122);border:1px #5f6368 solid;padding:0}.LGgmyb{bottom:0;left:0;opacity:0;position:absolute;right:0;top:0}.RpYYWb:not(.RDPZE) .LGgmyb{background-color:#3c4043}.kzYc3e:not(.RDPZE) .LGgmyb{background-color:#dadce0}.RpYYWb:hover .LGgmyb{opacity:0.04}.RpYYWb:focus .LGgmyb{opacity:0.12}.RpYYWb.u3bW4e:hover .LGgmyb{opacity:0.155}.kzYc3e:hover .LGgmyb{opacity:0.04}.kzYc3e:focus .LGgmyb{opacity:0.12}.kzYc3e.u3bW4e:hover .LGgmyb{opacity:0.155}.Qp3Dee{background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;transform:translate(-50%,-50%) scale(0);transition:opacity .2s ease,visibility 0s ease .2s,transform 0s ease .2s;transition:opacity .2s ease,visibility 0s ease .2s,-webkit-transform 0s ease .2s;top:0;visibility:hidden}.EijSib.qs41qe .Qp3Dee{opacity:1;transform:translate(-50%,-50%) scale(2.2);visibility:visible}.EijSib.qs41qe.M9Bg4d .Qp3Dee{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1),opacity .2s cubic-bezier(0,0,0.2,1)}.EijSib.j7nIZb .Qp3Dee{transform:translate(-50%,-50%) scale(2.2);visibility:visible}.RpYYWb .Qp3Dee{background-image:radial-gradient(circle farthest-side,rgba(60,64,67,0.102),rgba(60,64,67,0.102) 80%,rgba(60,64,67,0) 100%)}.kzYc3e .Qp3Dee{background-image:radial-gradient(circle farthest-side,rgba(218,220,224,0.102),rgba(218,220,224,0.102) 80%,rgba(218,220,224,0) 100%)}.f6aXTd{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;position:relative;margin:0 12px}.YcK5we{color:inherit;display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;fill:inherit;flex-shrink:0;margin:0 4px 0 -4px}.EijSib:not(.RDPZE).fy1E5c .YcK5we{color:#1a73e8;fill:#1a73e8}.kzYc3e:not(.RDPZE).fy1E5c .YcK5we{color:#8ab4f8;fill:#8ab4f8}.WUc8Ge.WUc8Ge{margin-right:-10px;width:28px;height:28px}.WUc8Ge:before{bottom:-10px;content:"";height:48px;left:-10px;position:absolute;right:-10px;top:-10px;width:48px}.f6aXTd .rag0{display:inline-block;margin:6px 4px}.hf2LYd{color:rgb(32,33,36);font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:2.75rem;font-size:2.25rem;letter-spacing:0;font-weight:400}.tl5cWb{color:rgb(32,33,36);font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:2.25rem;font-size:1.75rem;letter-spacing:0;font-weight:400}.FMcyT{color:rgb(32,33,36);font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.75rem;font-size:1.375rem;letter-spacing:0;font-weight:400}.Kqfayb{color:rgb(32,33,36);font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:500}.BgHQ3e{color:rgb(32,33,36);font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.xUvfQb{color:rgb(60,64,67);font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.0125em;font-weight:500}.w7mMgb{color:rgb(60,64,67);font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.XDCFvf{color:rgb(60,64,67);font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400}.FMzRdf{color:rgb(60,64,67);font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400}.MuGjgf{color:rgb(95,99,104);font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400}.qVzWGe{color:inherit;font-family:inherit;font-size:inherit;font-weight:inherit;letter-spacing:inherit;line-height:inherit}.QGK5hf{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:500}.jEt4Gf{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.mGD88b{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400}.eaF3Ie,.eaF3Ie:visited{color:rgb(25,103,210);cursor:pointer;text-decoration:none}.eaF3Ie:hover,.eaF3Ie:focus{outline:none;text-decoration:underline}.RMrItf{color:rgb(95,99,104)}.Vn3w8c{color:rgba(0,0,0,.38)}.Dcm1fd{color:rgb(217,48,37);font-style:italic}.VAPGpe{font-size:.1rem;height:.1rem;line-height:1;opacity:.001;overflow:hidden;position:absolute;width:.1rem}.K0lUWd{text-overflow:ellipsis;-o-text-overflow:ellipsis;-ms-text-overflow:ellipsis;overflow:hidden;white-space:nowrap;display:block}.sKKyEc{display:block;margin:-12px -12px}.pAlOFe{color:rgb(26,115,232);fill:rgb(26,115,232)}.Lzvjbf{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-flow:row nowrap}.XM8TV{-moz-box-flex:1;flex:1 0 4px}.ryQTbf{-moz-box-flex:1;flex:1 0 8px}.NHp4Tc{-moz-box-flex:1;flex:1 0 16px}.ft5Sbf{border:1px solid rgba(0,0,0,.12);border-radius:8px}.C4yF5e{border:1px solid rgba(0,0,0,.12);border-radius:4px}.EutHWe{-moz-box-align:center;align-items:center;display:-moz-box;display:flex}.LdvLn .snByac{text-overflow:ellipsis;-o-text-overflow:ellipsis;-ms-text-overflow:ellipsis;overflow:hidden;white-space:nowrap;text-align:left}.nmr34b .snByac{overflow:hidden}.nmr34b .Ce1Y1c,.k5SYqb .snByac{line-height:1.25rem}.YWEHbb{margin-left:8px}.PhlOZb{margin:0 -4px;padding:0 4px;font-style:italic}.xjQr1{height:16px;width:16px}.xjQr1 .GOJTSe{border-width:2px}.g4krrc.u3bW4e{outline:1px solid transparent}.wLnL5b{background-color:rgba(0,0,0,.12)!important}.oC328b{background-color:rgba(0,0,0,.24)!important}.C2NJgb{transition:background-color 0.28s 150ms}.C2NJgb>.DPvwYc{opacity:1;transition:opacity 0.28s 150ms}.wLnL5b.C2NJgb>.DPvwYc{opacity:0}.C9xz{display:inline-block;margin-bottom:.5rem;width:-moz-fit-content;width:fit-content}.szB9Tb,.szB9Tb:active,.szB9Tb:visited{color:inherit;text-decoration:none}.F4Rgre{max-width:100%}.aBlSgd{display:-moz-box;display:flex;margin-bottom:.5rem;margin-left:1rem;margin-right:1rem}.aBlSgd .rNj4oc{-moz-box-flex:1;flex-grow:1;width:0}.kg6ice{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.zZ8fDe{max-width:35rem}.qj5L0{border-bottom:.0625rem solid rgb(218,220,224);margin-bottom:.5rem;padding-bottom:1rem}.xhoYVc{padding-top:1rem}.jDlKLb{font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400;color:rgb(95,99,104);font-style:italic;margin-top:.625rem;text-align:center}.TH8fHb{margin-bottom:.875rem}.pjRund{-moz-box-orient:horizontal;-moz-box-direction:reverse;flex-direction:row-reverse}.pjRund .jDlKLb{margin-right:.625rem;margin-top:0;min-width:12.5rem;text-align:right}.Z3qXvc{margin:0 auto;max-width:47.5rem;padding:1.5rem 1.5rem}@media (max-width:30em){.Z3qXvc{width:auto;flex-direction:column;padding:0.5rem 0.5rem}}@media not all and (max-width:80.875em){.BdCNc{margin:1.5rem auto;width:-moz-calc(100% - 2*1.5rem);width:calc(100% - 2*1.5rem);max-width:47.5rem;position:relative}.GP1o5c{position:absolute;left:-14.625rem}}@media (max-width:80.875em){.GP1o5c{flex-shrink:0}.GP1o5c .asCVDb{margin-right:1.5rem}.BdCNc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;margin:1.5rem 1.5rem}.ihrflc{box-flex:1;flex-grow:1;max-width:47.5rem;min-width:0}}@media not all and (max-width:60rem){.smtc7c{display:none}}@media (max-width:60rem){.BdCNc{display:block;margin:1.5rem auto;padding:0 1.5rem;max-width:47.5rem;width:auto}.asCVDb{display:none}.A90zEf{display:block}}@media (max-width:48.75em){.pEwOBc{margin:0 -1.5rem}}@media (max-width:30em){.BdCNc{margin:0.5rem 0.5rem;padding:0}.pEwOBc{margin:0 -0.5rem}}.BdCNc.OOnEBd{position:static}.jeczbd:not(:empty)~*{display:none}.jeczbd:not(:empty){padding-bottom:0.5rem}.heSgkb{text-align:right}.uodSNb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;opacity:0.87}@media (max-width:40em){.aEqmgd{-moz-flex-wrap:wrap;flex-wrap:wrap}}.RpDEo{min-width:5.75rem}.yHjGtf{border-left:0.0625rem solid #e0e0e0;min-width:3.9375rem;padding:0 1rem;flex-shrink:0;text-decoration:none}.RpDEo{flex-shrink:0;text-decoration:none}.yHjGtf:focus{outline:none}.RpDEo:hover .J4BFhf,.RpDEo:focus .J4BFhf{color:#1a73e8;outline:none}.AXJKRe .J4BFhf{color:#9aa0a6}.GtqMq{cursor:default}.AsoHne{border-bottom:0.0625rem solid rgba(0,0,0,.87);display:inline-block;line-height:1;vertical-align:top;width:1.25rem}.ksaOtd{font-weight:500;color:rgba(0,0,0,.87)}.u7S8tc .DPvwYc{display:block}.UhYXkc{display:-ms-grid;display:grid}.u7S8tc+.E70Hue{pointer-events:none}.u7S8tc,.E70Hue{transition:opacity 0.28s cubic-bezier(0.4,0,0.2,1);grid-area:1/1}.u7S8tc{opacity:0;position:relative}.u7S8tc .WG5SSb{right:0;top:0}.ZnNi8e .E70Hue{opacity:0}.ZnNi8e .u7S8tc{opacity:1}.T0FFIe{font-size:0.875rem;font-weight:500;padding-left:1.5rem}.tfGBod.Yak70{border:none}.tfGBod:not(:first-child).kKn9Nc,.tfGBod.kKn9Nc+.tfGBod{border-top:none}.ubqkMe .jWCzBe .iobNdf,.J2ZeGc .jWCzBe .iobNdf,.svdjhb .jWCzBe .iobNdf{background-color:#bdc1c6}.D3ZbAb{flex-shrink:0;margin-right:1rem}.iobNdf{align-items:center;color:#fff;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:2.25rem;justify-content:center;margin-left:1.5rem;width:2.25rem}.FVAqmc .iobNdf{margin-left:0}.ubqkMe .kByKEb,.RyF19b .kByKEb,.J2ZeGc .kByKEb,.svdjhb .kByKEb{color:#5f6368}.ubqkMe .wCDkmf,.RyF19b .wCDkmf,.J2ZeGc .wCDkmf{font-style:italic}.RyF19b .wCDkmf,.RyF19b .iobNdf>.wVTR9d{color:#dd2c00}.kByKEb{width:100%}.tfGBod.xp2dJ{-moz-box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);list-style:none;max-width:-moz-calc(100% - (2*0.5rem));max-width:calc(100% - (2*0.5rem));width:17.5rem}.tfGBod.xp2dJ:before{-moz-box-shadow:none;box-shadow:none}.tfGBod.xp2dJ .a2rP{display:none}.tfGBod.tfGBod:not(.xp2dJ),.tfGBod.xp2dJ .jWCzBe,.tfGBod.xp2dJ .iobNdf{background-color:transparent}.tfGBod.J2ZeGc.xp2dJ,.tfGBod.ubqkMe.xp2dJ,.tfGBod.RyF19b.xp2dJ{background-color:#dadce0}.tfGBod.tfGBod.J2ZeGc.xp2dJ .iobNdf,.tfGBod.tfGBod.ubqkMe.xp2dJ .iobNdf{color:#3c4043;fill:#3c4043}.tfGBod.tfGBod.J2ZeGc.xp2dJ .xVnXCf *,.tfGBod.tfGBod.ubqkMe.xp2dJ .xVnXCf *,.tfGBod.tfGBod.RyF19b.xp2dJ .xVnXCf *{color:#3c4043}.tfGBod.xp2dJ .T3FW5d{display:none}.tfGBod.xp2dJ,.tfGBod.xp2dJ .jWCzBe{-moz-border-radius:0.5rem;border-radius:0.5rem;overflow:hidden}.tfGBod.xp2dJ .lio3ib{-moz-box-flex:1 1 auto;flex:1 1 auto}.tfGBod:not(.RyF19b).xp2dJ .jWCzBe *{color:white}.tfGBod.rZXyy:hover{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);border-radius:0.5rem;overflow:hidden}.tfGBod.rZXyy:not(.xp2dJ):hover .jWCzBe{background-color:white}.tfGBod.lXuxY.xp2dJ .jWCzBe{border-bottom:transparent}.tfGBod.lXuxY .jWCzBe .lio3ib{flex-basis:100%;flex-shrink:1;width:100%}.tfGBod.lXuxY .nZCyt{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.wvNVNd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row}.IMcm2d{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;margin-top:1rem}.bqKF7d,.vGGYOe{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:1;flex-grow:1;margin-left:0;min-width:0;overflow:hidden;text-overflow:ellipsis}.yVyYEc:not(:empty){margin-top:0.75rem}.rYHrHc{display:none}.a2rP .rYHrHc{display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;margin:-0.25rem 0}.KQqSid,.HSe5uf{box-flex:0;flex-grow:0;flex-shrink:0;margin-left:1rem}.O9YpHb:empty{display:none}.O9YpHb{border-top:0.0625rem solid #e0e0e0;box-sizing:border-box;flex-shrink:0;height:3.75rem;justify-content:space-between;padding:1rem 1.5rem}.mnp1de:not(:empty),.h3nrk:not(:empty){margin-top:1rem}.mnp1de{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;gap:1rem}.pSFXVb .LlHJB:not(:empty){margin-top:1.5rem}.uStMnd .bs9m7d:not(:empty){margin-top:1rem}.Mumuv{margin-bottom:1rem;margin-top:1rem}.FVAqmc .b9xlif{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:100%;position:absolute;right:0.5rem;top:0}.FVAqmc .b9xlif .ORmQmd{margin:0}.FVAqmc .bjejzf{padding-left:1.5rem;padding-right:-moz-calc(1rem + 48px);padding-right:calc(1rem + 48px)}.FVAqmc .bjejzf .lio3ib{-moz-box-flex:1 1 100%;flex:1 1 100%}.FVAqmc .jWCzBe .WZkEbf{font-size:0.875rem;font-weight:normal}.FVAqmc .IMcm2d{flex-direction:column}.FVAqmc .bqKF7d:not(:empty)+.KQqSid{margin-top:1rem}.FVAqmc .KQqSid{margin-left:0}.lio3ib{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:0 0 50%;flex:0 0 50%;flex-direction:column;min-width:0}.xVnXCf{height:100%;width:-moz-calc(100% - 4.75rem - 2.5rem - 1rem);width:calc(100% - 4.75rem - 2.5rem - 1rem)}.wCDkmf{box-sizing:border-box;color:rgba(0,0,0,.549);-moz-box-flex:0 0;flex:0 0;flex-basis:calc(30% - 1rem + 0.25rem);margin-left:1rem;min-width:0;padding-right:0.25rem;margin-right:-0.25rem;text-align:right}.nZCyt{color:rgba(0,0,0,.549);-moz-box-flex:0 0;flex:0 0;flex-basis:calc(20% - 1rem);margin-left:1rem;min-width:0}@media (max-width:30em){.jWCzBe .wCDkmf,.jWCzBe .nZCyt{display:none}.jWCzBe .lio3ib{-moz-box-flex:0 0 100%;flex:0 0 100%}}@media not all and (max-width:30em){.jWCzBe .WZkEbf{display:none}}.WZkEbf:not(:empty){margin-top:0.25rem}.WyjGac{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:0;flex-grow:0;flex-shrink:0;justify-content:center;margin:0 0.5rem;width:2.5rem}.zIKt9b .lGm3nb .JRtysb{color:transparent;fill:transparent}.jWCzBe:hover .lGm3nb .I12f0b,.jWCzBe:focus .lGm3nb .I12f0b,.xVnXCf:focus+.WyjGac .I12f0b,.lGm3nb .I12f0b.iWO5td,.lGm3nb .I12f0b:focus{color:#5f6368;fill:#5f6368}.yPNvqb{color:transparent}.yPNvqb .Vk3rb .DPvwYc{color:rgba(0,0,0,.549)}.jWCzBe:hover .yPNvqb,.jWCzBe:focus .yPNvqb{color:#444}.DzHQo{position:relative}.GfOiTd,.b5T4ud{color:rgba(0,0,0,.549);display:-moz-box;display:flex;padding:1rem 1.5rem}.eSRRRc .GfOiTd{display:none}.eSRRRc .Xzp3fc{min-height:3.75rem}.eSRRRc .kKn9Nc{background-color:transparent;position:relative;visibility:visible}.eSRRRc .kKn9Nc *{visibility:hidden}.eSRRRc .kKn9Nc:before{background-color:rgb(241,243,244);border-radius:.5rem;bottom:0;box-shadow:none;content:"";left:0;position:absolute;right:0;top:0;z-index:0}.eSRRRc .Xzp3fc:after{content:"";display:block;height:3.75rem;margin-bottom:-3.75rem;width:100%}.eSRRRc .a2rP{display:none}.eSRRRc .tfGBod.Oan9Gc,.eSRRRc .tfGBod.Oan9Gc+.tfGBod{border-top:none;margin-top:0}.GfOiTd,.b5T4ud{-moz-box-align:center;align-items:center;-moz-box-sizing:border-box;box-sizing:border-box;height:3.75rem;z-index:0}.Mvr5Ef{display:-moz-box;display:flex;-moz-box-pack:center;justify-content:center;min-height:.5rem}.nZ34k{margin-bottom:.25rem;margin-top:.25rem}.nZ34k:not(:disabled){color:#5f6368}.nZ34k:not(:disabled):hover{color:#5f6368}.nZ34k:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.nZ34k:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:#5f6368}.iBZDFb{top:-2.5px;left:0;position:absolute;right:0;width:100%}.fwcY1d{cursor:pointer;padding:0 1.5rem}.ovsVve[aria-expanded="true"] .fwcY1d{margin-bottom:1rem}@media (max-width:30em){.ovsVve[aria-expanded="true"] .fwcY1d{margin-bottom:0.5rem}.fwcY1d{padding:0.5rem 1rem}}.vU3YFf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-right:0.75rem}.ovsVve.Aopndd .fwcY1d{margin-bottom:0;padding:0.5rem 1rem}.ovsVve.Aopndd .JQIfHf{padding:0.5rem 1rem}.KmLLod:hover{-moz-border-radius:0.5rem;border-radius:0.5rem}.KmLLod:hover .uO32ac{border-bottom:none}.FpfvHe>.kKn9Nc{background-color:transparent;position:relative;visibility:visible}.FpfvHe>.kKn9Nc *{visibility:hidden}.FpfvHe>.kKn9Nc:before{background-color:#f1f3f4;-moz-border-radius:0.5rem;border-radius:0.5rem;bottom:0;-moz-box-shadow:none;box-shadow:none;content:"";left:0;position:absolute;right:0;top:0;z-index:0}.qdhuXb .FpfvHe:after{content:"";display:block;height:3.75rem;margin-bottom:-3.75rem;width:100%}.jHgkif.YwNp1:not(.xp2dJ){-moz-border-radius:0.5rem;border-radius:0.5rem;overflow:hidden}.jHgkif.YwNp1.xp2dJ{-moz-box-shadow:none;box-shadow:none}.jHgkif.xp2dJ .O1l69{-moz-border-radius:0.5rem;border-radius:0.5rem}.FpfvHe .jHgkif:not(.xp2dJ) .O1l69{background-color:transparent}.jHgkif.xp2dJ .O1l69 *{color:white}.jHgkif.xp2dJ .ClSQxf{display:none}.jHgkif.xp2dJ{-moz-box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);list-style:none;max-width:-moz-calc(100% - (2*0.5rem));max-width:calc(100% - (2*0.5rem));width:17.5rem}@media (max-width:40em){.qdhuXb .jHgkif:not(.xp2dJ) .zq2w8b{display:none}}.FpfvHe>.kKn9Nc .zq2w8b,.jHgkif.xp2dJ .zq2w8b{display:none}.jHgkif.xp2dJ{z-index:1100}.jHgkif.xp2dJ .O1l69{position:relative}.jHgkif.xp2dJ .O1l69:before{background:white;border:0.0625rem solid #e0e0e0;-moz-border-radius:0.5rem;border-radius:0.5rem;border-top:none;-moz-box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);content:"";position:absolute}.jHgkif.xp2dJ .O1l69:after{background:white;border:0.0625rem solid #e0e0e0;-moz-border-radius:0.5rem;border-radius:0.5rem;border-top:none;-moz-box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);content:"";position:absolute}.jHgkif.xp2dJ .O1l69:before{bottom:-0.5rem;left:0.5rem;right:-0.5rem;top:0.5rem;z-index:-1}.jHgkif.xp2dJ .O1l69:after{box-shadow:0 4px 4px 0 rgba(60,64,67,.3),0 8px 12px 6px rgba(60,64,67,.15);bottom:-1rem;left:1rem;right:-1rem;top:1rem;z-index:-2}.JBMs6{align-items:center;-moz-border-radius:0.5rem 0.5rem 0 0;border-radius:0.5rem 0.5rem 0 0;box-sizing:border-box;color:#fff;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;justify-content:space-between;padding:1.5rem}.jHgkif.xp2dJ .JBMs6.uO32ac{border-bottom:none}@media (max-width:40em){.qdhuXb .jHgkif .JBMs6.uO32ac{border-bottom:none}}.ClSQxf{margin-right:-1rem}.xUYklb{margin:-1rem 0 -1rem -1.5rem;padding:1rem 0 1rem 1.5rem;text-decoration:none;width:100%}.jHgkif .ovsVve .fwcY1d{box-sizing:border-box;height:3.75rem;padding:1.5rem}.jHgkif .ovsVve[aria-expanded="true"] .fwcY1d{margin-bottom:0}.jHgkif .ovsVve[aria-expanded="true"]{background-color:transparent;padding:0}.JZINBb{border-bottom:0.0625rem solid #e0e0e0;border-width:0.125rem;margin-top:2.5rem}.Ju84Lc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;margin:8.4375rem 0 1.5rem}.bqfGyf{height:7.1875rem}.m5Cxw{margin-bottom:0.5rem;text-align:center}.z4rkrb{margin:0 auto 2rem;max-width:21.875rem;text-align:center}.k2wCFc{flex-direction:row}.tCD5Mc{flex-shrink:1;padding:1.5rem 1.5rem 0;margin:1rem 1.5rem;width:24rem}.tCD5Mc h1{margin-bottom:1rem}.tCD5Mc p{margin-bottom:1.5rem;margin-top:0}.QWwQ3c{margin-bottom:1rem;justify-content:flex-end;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:wrap;flex-wrap:wrap}.QWwQ3c>.QRiHXd{justify-content:flex-end;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:wrap;flex-wrap:wrap}.QWwQ3c .ZSrdFd,.QWwQ3c .uArJ5e{margin-bottom:0.5rem;margin-left:1rem;margin-right:0;text-decoration:none}.r8WYMb{margin-bottom:0.5rem;margin-top:-14px}.FHIL6b{margin-bottom:1rem}.xd70xe:not(:empty){margin-bottom:1rem;word-wrap:break-word}.V8apv{background-color:#f8f9fa;-moz-border-radius:0.5rem;border-radius:0.5rem}.GOm7re{-moz-flex-wrap:wrap;flex-wrap:wrap}.GOm7re>*:not(:empty){margin-bottom:1rem}.GOm7re .oxacD.oxacD{margin-top:0}.X4kONd{margin-bottom:1rem;width:100%}.ITx4Gf{-moz-box-ordinal-group:1;order:1}.r1i1xd{margin-right:1rem;max-width:25rem;-moz-box-ordinal-group:2;order:2}.GAU0yc{-moz-box-ordinal-group:3;order:3}.Im5hIb{text-align:center}.e6es3,.XfQwid{display:none}.JZgRpf .e6es3,.q163ye .XfQwid{display:block}.jlVFDe{margin-bottom:1rem;line-height:1}.eaNNh{display:inline-block;margin:0 .5rem}.HMTQQd{margin:-.625rem -.5rem;opacity:.54}.MGdB9c{margin-bottom:1.5rem}.ZQXs7e.eiJHkc{border-bottom-right-radius:0;border-top-right-radius:0;margin-right:.0625rem}@media not all and (max-width:40rem){.ZQXs7e.qs9Ooe{border-bottom-right-radius:0;border-top-right-radius:0;margin-right:.0625rem}}.nNUyy{align-self:stretch;border-bottom-left-radius:0;border-top-left-radius:0;display:-moz-box;display:flex;-moz-box-pack:center;justify-content:center;min-width:2.125rem}.A8QgL.A8QgL{margin-left:.5rem}.nNUyy .Fxmcue{padding:0 .25rem}.nNUyy .snByac{-moz-box-align:center;align-items:center;display:-moz-box;display:flex}.wMkDgf{font-style:italic;flex-shrink:0;margin-right:1rem}@media not all and (max-width:40em){.S5j4t{margin-right:0.5rem}}.HvC6Tb{display:-moz-box;display:flex;overflow:hidden}.e0prFf{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.75rem;font-size:1.375rem;letter-spacing:0;font-weight:400;color:rgb(95,99,104);-moz-box-flex:1;flex-grow:1;min-width:0;padding:.25rem;padding-left:.75rem}.XpCIle{height:2.25rem;width:2.25rem}.efOAcd{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;flex-shrink:0}.wyl3j{z-index:3000}.UsVAVe{border-color:rgb(232,234,237);border-radius:50%;border-style:solid;border-width:.0625rem;height:3rem;margin:.625rem .5rem;width:3rem}.C3VsHd{height:1.5rem;width:1.5rem}.gGXFW{max-width:980px;width:100%}.mstpre.z80M1.FeRvI{padding-left:0}.jwVv6b{margin-left:8px}.pFwdNe{max-height:13.75rem;overflow:auto;width:100%}.pFwdNe .LoI3h{border-radius:.4375rem}.pFwdNe .LoI3h.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:44px}.pFwdNe .LoI3h.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.pFwdNe .LoI3h.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:60px}.vI34tf{display:inline-block;height:100%;width:100%}.gCiH5e{padding-top:.625rem;text-align:center;width:100%}.VlVMqe{height:4.0625rem;margin-bottom:.625rem}.lLyPQd{margin-bottom:2.8125rem;margin-top:0}.v58QK{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;margin-bottom:.3125rem}.qplEpd{font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400;font-style:italic;color:rgb(95,99,104);margin-bottom:1.25rem}.Di7vwd{width:44px;height:44px;padding:11px;font-size:22px;background:#fff;border-radius:1.5625rem;margin-right:.25rem;opacity:0;padding:.5rem 0 0 .25rem;position:absolute;right:0;top:-.125rem}.Di7vwd svg,.Di7vwd img{width:22px;height:22px}.LoI3h:active .Di7vwd,.Di7vwd:active{background:rgb(218,220,224)}.LoI3h:hover .Di7vwd,.LoI3h:focus .Di7vwd,.Di7vwd:hover,.Di7vwd:focus{color:rgb(95,99,104);display:inline-block;-moz-box-pack:center;justify-content:center;pointer-events:auto;opacity:1}@media (max-width:30rem){.Di7vwd{opacity:1}}.KkCUjb{height:2.5rem;min-width:12.5rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::before,.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-mWPk3d .VfPpkd-fmcmS-OyKIhb::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-mWPk3d .VfPpkd-fmcmS-OyKIhb::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-fmcmS-OyKIhb::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-fmcmS-OyKIhb::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-fmcmS-OyKIhb::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::before,.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::after{top:-50%;left:-50%;width:200%;height:200%}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-mWPk3d .VfPpkd-fmcmS-OyKIhb::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-fmcmS-OyKIhb{position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}.VfPpkd-fmcmS-yrriRe{border-top-left-radius:4px;border-top-left-radius:var(--mdc-shape-small,4px);border-top-right-radius:4px;border-top-right-radius:var(--mdc-shape-small,4px);border-bottom-right-radius:0;border-bottom-left-radius:0;display:-moz-inline-box;display:inline-flex;-moz-box-align:baseline;align-items:baseline;padding:0 16px;position:relative;-moz-box-sizing:border-box;box-sizing:border-box;overflow:hidden;will-change:opacity,transform,color}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgba(0,0,0,.6)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgba(0,0,0,.87)}@media all{.mdc-text-field:not(.mdc-text-field--disabled) .mdc-text-field__input::-moz-placeholder{color:rgba(0,0,0,.54)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(0,0,0,.54)}}@media all{.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(0,0,0,.54)}}.VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-wGMbrd{caret-color:#6200ee;caret-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgba(0,0,0,.6)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(0,0,0,.6)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgba(0,0,0,.54)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(0,0,0,.54)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgba(0,0,0,.6)}.VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(0,0,0,.6)}.VfPpkd-fmcmS-yrriRe .VfPpkd-NLUYnc-V67aGc{top:50%;transform:translateY(-50%);pointer-events:none}.VfPpkd-fmcmS-wGMbrd{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);height:28px;transition:opacity .15s 0ms cubic-bezier(.4,0,.2,1);width:100%;min-width:0;border:none;border-radius:0;background:none;-moz-appearance:none;appearance:none;padding:0}.VfPpkd-fmcmS-wGMbrd::-ms-clear{display:none}.VfPpkd-fmcmS-wGMbrd::-webkit-calendar-picker-indicator{display:none}.VfPpkd-fmcmS-wGMbrd:focus{outline:none}.VfPpkd-fmcmS-wGMbrd:invalid{box-shadow:none}@media all{.mdc-text-field__input::-moz-placeholder{-moz-transition:opacity 67ms 0ms cubic-bezier(.4,0,.2,1);transition:opacity 67ms 0ms cubic-bezier(.4,0,.2,1);opacity:0}.VfPpkd-fmcmS-wGMbrd::placeholder{transition:opacity 67ms 0ms cubic-bezier(.4,0,.2,1);opacity:0}}@media all{.VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{-ms-transition:opacity 67ms 0ms cubic-bezier(.4,0,.2,1);transition:opacity 67ms 0ms cubic-bezier(.4,0,.2,1);opacity:0}}@media all{.mdc-text-field--no-label .mdc-text-field__input::-moz-placeholder, .mdc-text-field--focused .mdc-text-field__input::-moz-placeholder{transition-delay:40ms;transition-duration:.11s;opacity:1}.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc .VfPpkd-fmcmS-wGMbrd::placeholder,.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd::placeholder{transition-delay:40ms;transition-duration:.11s;opacity:1}}@media all{.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder,.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{transition-delay:40ms;transition-duration:.11s;opacity:1}}.VfPpkd-fmcmS-MvKemf{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);height:28px;transition:opacity .15s 0ms cubic-bezier(.4,0,.2,1);opacity:0;white-space:nowrap}.VfPpkd-fmcmS-yrriRe-OWXEXe-V67aGc-NLUYnc .VfPpkd-fmcmS-MvKemf,.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc .VfPpkd-fmcmS-MvKemf{opacity:1}@supports (-webkit-hyphens:none){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-MvKemf{-moz-box-align:center;align-items:center;align-self:center;display:-moz-inline-box;display:inline-flex;height:100%}}.VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{padding-left:0;padding-right:2px}[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c[dir=rtl]{padding-left:2px;padding-right:0}.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{padding-left:0;padding-right:12px}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c[dir=rtl]{padding-left:12px;padding-right:0}.VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{padding-left:12px;padding-right:0}[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB,.VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB[dir=rtl]{padding-left:0;padding-right:12px}.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{padding-left:2px;padding-right:0}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB,.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB[dir=rtl]{padding-left:0;padding-right:2px}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be{height:56px}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::before,.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb::after{background-color:rgba(0,0,0,.87);background-color:var(--mdc-ripple-color,rgba(0,0,0,.87))}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be:hover .VfPpkd-fmcmS-OyKIhb::before,.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-fmcmS-OyKIhb::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-fmcmS-OyKIhb::before,.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-fmcmS-OyKIhb::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be::before{display:inline-block;width:0;height:40px;content:"";vertical-align:0}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me){background-color:whitesmoke}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(0,0,0,.42)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(0,0,0,.87)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:#6200ee;border-bottom-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{left:16px;right:auto}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc,.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:16px}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-106%) scale(.75)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc .VfPpkd-fmcmS-wGMbrd{height:100%}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc .VfPpkd-NLUYnc-V67aGc{display:none}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc::before{display:none}@supports (-webkit-hyphens:none){.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc .VfPpkd-fmcmS-MvKemf{-moz-box-align:center;align-items:center;align-self:center;display:-moz-inline-box;display:inline-flex;height:100%}}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc{height:56px;overflow:visible}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-37.25px) scale(1)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:.75rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-34.75px) scale(.75)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:1rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-text-field-outlined .25s 1}@keyframes mdc-floating-label-shake-float-above-text-field-outlined{0%{transform:translateX(0) translateY(-34.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(4%) translateY(-34.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(-4%) translateY(-34.75px) scale(.75)}100%{transform:translateX(0) translateY(-34.75px) scale(.75)}}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-wGMbrd{height:100%}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(0,0,0,.38)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(0,0,0,.87)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-MpmGFe{border-color:#6200ee;border-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb{border-top-left-radius:4px;border-top-left-radius:var(--mdc-shape-small,4px);border-top-right-radius:0;border-bottom-right-radius:0;border-bottom-left-radius:4px;border-bottom-left-radius:var(--mdc-shape-small,4px)}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb[dir=rtl]{border-top-left-radius:0;border-top-right-radius:4px;border-top-right-radius:var(--mdc-shape-small,4px);border-bottom-right-radius:4px;border-bottom-right-radius:var(--mdc-shape-small,4px);border-bottom-left-radius:0}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb{width:max(12px,var(--mdc-shape-small,4px))}}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd{max-width:calc(100% - max(12px, var(--mdc-shape-small, 4px))*2)}}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-top-left-radius:0;border-top-right-radius:4px;border-top-right-radius:var(--mdc-shape-small,4px);border-bottom-right-radius:4px;border-bottom-right-radius:var(--mdc-shape-small,4px);border-bottom-left-radius:0}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe[dir=rtl]{border-top-left-radius:4px;border-top-left-radius:var(--mdc-shape-small,4px);border-top-right-radius:0;border-bottom-right-radius:0;border-bottom-left-radius:4px;border-bottom-left-radius:var(--mdc-shape-small,4px)}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc{padding-left:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc{padding-right:max(16px,var(--mdc-shape-small,4px))}}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc{padding-left:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc{padding-right:max(16px,var(--mdc-shape-small,4px))}}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c{padding-left:0}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c{padding-right:max(16px,var(--mdc-shape-small,4px))}}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c[dir=rtl]{padding-right:0}@supports (top:max(0%)){[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c[dir=rtl]{padding-left:max(16px,var(--mdc-shape-small,4px))}}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c{padding-right:0}@supports (top:max(0%)){.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c{padding-left:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c[dir=rtl]{padding-left:0}@supports (top:max(0%)){[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c[dir=rtl]{padding-right:max(16px,calc(var(--mdc-shape-small, 4px) + 4px))}}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c{padding-left:0;padding-right:0}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd{padding-top:1px}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-OyKIhb::before,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-OyKIhb::after{background-color:transparent;background-color:var(--mdc-ripple-color,transparent)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc{left:4px;right:auto}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:4px}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-wGMbrd{display:-moz-box;display:flex;border:none!important;background-color:transparent}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e{z-index:1}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od{-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-align:center;align-items:center;width:auto;height:auto;padding:0;transition:none}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od .VfPpkd-NLUYnc-V67aGc{top:19px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od .VfPpkd-NLUYnc-V67aGc:not(.VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe){transform:none}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od .VfPpkd-fmcmS-wGMbrd{-moz-box-flex:1;flex-grow:1;height:auto;min-height:1.5rem;overflow-x:hidden;overflow-y:auto;-moz-box-sizing:border-box;box-sizing:border-box;resize:none;padding:0 16px;line-height:1.5rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be::before{display:none}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-10.25px) scale(.75)}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-textarea-filled .25s 1}@keyframes mdc-floating-label-shake-float-above-textarea-filled{0%{transform:translateX(0) translateY(-10.25px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(4%) translateY(-10.25px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(-4%) translateY(-10.25px) scale(.75)}100%{transform:translateX(0) translateY(-10.25px) scale(.75)}}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-wGMbrd{margin-top:23px;margin-bottom:9px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be.VfPpkd-fmcmS-yrriRe-OWXEXe-di8rgd-V67aGc .VfPpkd-fmcmS-wGMbrd{margin-top:16px;margin-bottom:16px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd{padding-top:0}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-27.25px) scale(1)}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:.75rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-24.75px) scale(.75)}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:1rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-textarea-outlined .25s 1}@keyframes mdc-floating-label-shake-float-above-textarea-outlined{0%{transform:translateX(0) translateY(-24.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(4%) translateY(-24.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(-4%) translateY(-24.75px) scale(.75)}100%{transform:translateX(0) translateY(-24.75px) scale(.75)}}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-wGMbrd{margin-top:16px;margin-bottom:16px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc{top:18px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-k4Qmrd-gmhCAd .VfPpkd-fmcmS-wGMbrd{margin-bottom:2px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-k4Qmrd-gmhCAd .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{align-self:flex-end;padding:0 16px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-k4Qmrd-gmhCAd .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd::after{display:inline-block;width:0;height:16px;content:"";vertical-align:-16px}.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-k4Qmrd-gmhCAd .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd::before{display:none}.VfPpkd-fmcmS-kHQaff{align-self:stretch;display:-moz-inline-box;display:inline-flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-flex:1;flex-grow:1;max-height:100%;max-width:100%;min-height:56px;min-width:-moz-fit-content;min-width:fit-content;min-width:-moz-available;min-width:-webkit-fill-available;overflow:hidden;resize:both}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-kHQaff{transform:translateY(-1px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-wGMbrd,.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{transform:translateY(1px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff{transform:translateX(-1px) translateY(-1px)}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff[dir=rtl]{transform:translateX(1px) translateY(-1px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-wGMbrd,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{transform:translateX(1px) translateY(1px)}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-wGMbrd,[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-wGMbrd[dir=rtl],.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-fmcmS-kHQaff .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd[dir=rtl]{transform:translateX(-1px) translateY(1px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c{padding-left:0;padding-right:16px}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c[dir=rtl]{padding-left:16px;padding-right:0}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{max-width:calc(100% - 48px);left:48px;right:auto}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:48px}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:calc(133.3333333333% - 85.3333333333px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc{left:36px;right:auto}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc[dir=rtl]{left:auto;right:36px}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc :not(.VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd) .VfPpkd-NSFCdd-Ra9xwd{max-width:calc(100% - 60px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-37.25px) translateX(-32px) scale(1)}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe[dir=rtl]{transform:translateY(-37.25px) translateX(32px) scale(1)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:.75rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-34.75px) translateX(-32px) scale(.75)}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe[dir=rtl],.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe[dir=rtl]{transform:translateY(-34.75px) translateX(32px) scale(.75)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:1rem}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-text-field-outlined-leading-icon .25s 1}@keyframes mdc-floating-label-shake-float-above-text-field-outlined-leading-icon{0%{transform:translateX(-32px) translateY(-34.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(calc(4% - 32px)) translateY(-34.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(calc(-4% - 32px)) translateY(-34.75px) scale(.75)}100%{transform:translateX(-32px) translateY(-34.75px) scale(.75)}}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc[dir=rtl] .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-text-field-outlined-leading-icon .25s 1}@keyframes mdc-floating-label-shake-float-above-text-field-outlined-leading-icon-rtl{0%{transform:translateX(32px) translateY(-34.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(calc(4% + 32px)) translateY(-34.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(calc(-4% + 32px)) translateY(-34.75px) scale(.75)}100%{transform:translateX(32px) translateY(-34.75px) scale(.75)}}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c{padding-left:16px;padding-right:0}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c,.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c[dir=rtl]{padding-left:0;padding-right:16px}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{max-width:calc(100% - 64px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:calc(133.3333333333% - 85.3333333333px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc :not(.VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd) .VfPpkd-NSFCdd-Ra9xwd{max-width:calc(100% - 60px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c{padding-left:0;padding-right:0}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{max-width:calc(100% - 96px)}.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:calc(133.3333333333% - 128px)}.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc{display:-moz-box;display:flex;-moz-box-pack:justify;justify-content:space-between;-moz-box-sizing:border-box;box-sizing:border-box}.VfPpkd-fmcmS-yrriRe+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc{padding-right:16px;padding-left:16px}.VfPpkd-I9GLp-yrriRe>.VfPpkd-fmcmS-yrriRe+label{align-self:flex-start}.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgba(98,0,238,.87)}.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-MpmGFe{border-width:2px}.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS:not(.VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb){opacity:1}.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc .VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd{padding-top:2px}.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe.VfPpkd-fmcmS-yrriRe-OWXEXe-INsAgc.VfPpkd-fmcmS-yrriRe-OWXEXe-B7I4Od .VfPpkd-NSFCdd-i5vt6e-OWXEXe-NSFCdd .VfPpkd-NSFCdd-Ra9xwd{padding-top:0}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:#b00020;border-bottom-color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:#b00020;border-bottom-color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:#b00020;color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:#b00020;color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:#b00020;caret-color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:#b00020;color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:#b00020;border-bottom-color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:#b00020;border-color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:#b00020;border-color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NSFCdd-MpmGFe{border-color:#b00020;border-color:var(--mdc-theme-error,#b00020)}.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{opacity:1}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me{pointer-events:none}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(0,0,0,.38)}@media all{.mdc-text-field--disabled .mdc-text-field__input::-moz-placeholder{color:rgba(0,0,0,.38)}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(0,0,0,.38)}}@media all{.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(0,0,0,.38)}}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(0,0,0,.38)}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(0,0,0,.3)}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(0,0,0,.38)}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(0,0,0,.06)}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(0,0,0,.06)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.mdc-text-field--disabled .mdc-text-field__input::-moz-placeholder{color:GrayText}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:GrayText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:GrayText}}@media screen and (forced-colors:active){.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{background-color:Window}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{z-index:1}}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{cursor:default}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be{background-color:#fafafa}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me.VfPpkd-fmcmS-yrriRe-OWXEXe-MFS4be .VfPpkd-fmcmS-OyKIhb{display:none}.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{pointer-events:auto}.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-wGMbrd{text-align:right}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-wGMbrd,.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-wGMbrd[dir=rtl]{text-align:left}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-wGMbrd,[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-MvKemf,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-wGMbrd,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-MvKemf{direction:ltr}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{padding-left:0;padding-right:2px}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{padding-left:12px;padding-right:0}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{-moz-box-ordinal-group:2;order:1}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{-moz-box-ordinal-group:3;order:2}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-wGMbrd,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-wGMbrd{-moz-box-ordinal-group:4;order:3}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{-moz-box-ordinal-group:5;order:4}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS[dir=rtl] .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{-moz-box-ordinal-group:6;order:5}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-wGMbrd,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd[dir=rtl] .VfPpkd-fmcmS-wGMbrd{text-align:right}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{padding-right:12px}[dir=rtl] .VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB,.VfPpkd-fmcmS-yrriRe-OWXEXe-i3jM8c-fmcmS.VfPpkd-fmcmS-yrriRe-OWXEXe-CpWD9d-KW5YQd[dir=rtl] .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{padding-left:2px}.VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit);display:block;margin-top:0;line-height:normal;margin:0;opacity:0;will-change:opacity;transition:opacity .15s 0ms cubic-bezier(.4,0,.2,1)}.VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS::before{display:inline-block;width:0;height:16px;content:"";vertical-align:0}.VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS-OWXEXe-zvnfze{transition:none;opacity:1;will-change:auto}.VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit);display:block;margin-top:0;line-height:normal;margin-left:auto;margin-right:0;padding-left:16px;padding-right:0;white-space:nowrap}.VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd::before{display:inline-block;width:0;height:16px;content:"";vertical-align:0}[dir=rtl] .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd[dir=rtl]{margin-left:0;margin-right:auto}[dir=rtl] .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd[dir=rtl]{padding-left:0;padding-right:16px}.VfPpkd-fmcmS-TvZj5c{align-self:center;cursor:pointer}.VfPpkd-fmcmS-TvZj5c:not([tabindex]),.VfPpkd-fmcmS-TvZj5c[tabindex="-1"]{cursor:default;pointer-events:none}.VfPpkd-fmcmS-TvZj5c svg{display:block}.VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{margin-left:16px;margin-right:8px}[dir=rtl] .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc[dir=rtl]{margin-left:8px;margin-right:16px}.VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{padding:12px;margin-left:0;margin-right:0}[dir=rtl] .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg,.VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg[dir=rtl]{margin-left:0;margin-right:0}.WmnPA+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS,.WmnPA+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400;line-height:.875rem}.WmnPA .VfPpkd-NLUYnc-V67aGc{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;line-height:1.15rem}.WmnPA .VfPpkd-fmcmS-wGMbrd{font-family:Roboto,Arial,sans-serif;font-size:1rem;letter-spacing:.00625em;font-weight:400}.WmnPA:hover .VfPpkd-fmcmS-OyKIhb::before,.WmnPA.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-fmcmS-OyKIhb::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.WmnPA.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-fmcmS-OyKIhb::before,.WmnPA:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-fmcmS-OyKIhb::before{transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.WmnPA .VfPpkd-fmcmS-OyKIhb::before,.WmnPA .VfPpkd-fmcmS-OyKIhb::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(95,99,104)}.WmnPA .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(25,103,210)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(60,64,67)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me){background-color:rgb(241,243,244)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(95,99,104)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(95,99,104)}.WmnPA:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(32,33,36)}.WmnPA:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(32,33,36)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(95,99,104)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(25,103,210)}@media all{.GmTextFieldBox:not(.mdc-text-field--disabled) .mdc-text-field__input::-moz-placeholder{color:rgb(95,99,104)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(95,99,104)}}@media all{.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(95,99,104)}}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(95,99,104)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(95,99,104)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(95,99,104)}.WmnPA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(95,99,104)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(60,64,67,.38)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me{background-color:rgba(95,99,104,.04)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(95,99,104,.38)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(95,99,104,.38)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(60,64,67,.38)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgba(95,99,104,.38)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(60,64,67,.38)}@media all{.GmTextFieldBox.mdc-text-field--disabled .mdc-text-field__input::-moz-placeholder{color:rgba(60,64,67,.38)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(60,64,67,.38)}}@media all{.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(60,64,67,.38)}}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(60,64,67,.38)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(25,103,210)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(197,34,31)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(197,34,31)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(217,48,37)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(197,34,31)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(197,34,31)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(165,14,14)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(165,14,14)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(165,14,14)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(165,14,14)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(25,103,210)}.WmnPA.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(197,34,31)}.cfWmIb+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS,.cfWmIb+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400;line-height:.875rem}.cfWmIb .VfPpkd-NLUYnc-V67aGc{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;line-height:1.15rem}.cfWmIb .VfPpkd-fmcmS-wGMbrd{font-family:Roboto,Arial,sans-serif;font-size:1rem;letter-spacing:.00625em;font-weight:400}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(60,64,67);color:var(--gm-outlinedtextfield-ink-color,rgb(60,64,67))}.cfWmIb .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(26,115,232);caret-color:var(--gm-outlinedtextfield-caret-color,rgb(26,115,232))}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-helper-text-color,rgb(95,99,104))}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(95,99,104)}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-label-color,rgb(95,99,104))}.cfWmIb:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(32,33,36)}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(128,134,139);border-color:var(--gm-outlinedtextfield-outline-color,rgb(128,134,139))}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(32,33,36)}@media all{.GmTextFieldOutlined:not(.mdc-text-field--disabled) .mdc-text-field__input::-moz-placeholder{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-placeholder-color,rgb(95,99,104))}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-placeholder-color,rgb(95,99,104))}}@media all{.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-placeholder-color,rgb(95,99,104))}}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-prefix-color,rgb(95,99,104))}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-suffix-color,rgb(95,99,104))}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(95,99,104)}.cfWmIb:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(95,99,104)}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-ink-color--disabled,rgba(95,99,104,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(60,64,67,.12);border-color:var(--gm-outlinedtextfield-outline-color--disabled,rgba(60,64,67,.12))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-label-color--disabled,rgba(95,99,104,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(95,99,104,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(95,99,104,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-helper-text-color--disabled,rgba(95,99,104,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-character-counter-color--disabled,rgba(95,99,104,.38))}@media all{.GmTextFieldOutlined.mdc-text-field--disabled .mdc-text-field__input::-moz-placeholder{color:rgba(60,64,67,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(60,64,67,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(60,64,67,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(60,64,67,.38))}}@media all{.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(60,64,67,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(60,64,67,.38))}}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-prefix-color--disabled,rgba(95,99,104,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-suffix-color--disabled,rgba(95,99,104,.38))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(26,115,232);border-color:var(--gm-outlinedtextfield-outline-color--stateful,rgb(26,115,232))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(26,115,232);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(26,115,232))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(217,48,37);caret-color:var(--gm-outlinedtextfield-caret-color--error,rgb(217,48,37))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(217,48,37);color:var(--gm-outlinedtextfield-helper-text-color--error,rgb(217,48,37))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(165,14,14)}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(165,14,14)}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(165,14,14)}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(165,14,14)}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(217,48,37);border-color:var(--gm-outlinedtextfield-outline-color--error,rgb(217,48,37))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(217,48,37);color:var(--gm-outlinedtextfield-icon-color--error,rgb(217,48,37))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(217,48,37);border-color:var(--gm-outlinedtextfield-outline-color--error-stateful,rgb(217,48,37))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(26,115,232);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(26,115,232))}.cfWmIb.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(217,48,37);color:var(--gm-outlinedtextfield-label-color--error,rgb(217,48,37))}.cfWmIb .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:1rem}.cfWmIb .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:.75rem}.Tj45d{position:relative}.ncIyJc{position:absolute;overflow:hidden;left:-1px;top:auto;width:1px;height:1px}.Ufn6O{display:-moz-inline-box;display:inline-flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;position:relative}.Ufn6O[hidden]{display:none}.xlHPle{display:-moz-inline-box;display:inline-flex;position:relative}.xlHPle[hidden]{display:none}.xlHPle .UMrnmb-lP5Lpb-yrriRe,.xlHPle .UMrnmb-fdMfRe{width:inherit}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px}[dir=rtl] .xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.xlHPle .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:8px}[dir=rtl] .xlHPle .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc,.xlHPle .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:8px;margin-right:0}.xlHPle .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:48px;padding-right:16px}[dir=rtl] .xlHPle .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b,.xlHPle .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:48px}.xlHPle .VfPpkd-xl07Ob-XxIAqe-OWXEXe-uxVfW-FNFY6c-uFfGwd{border-top-left-radius:0;border-top-right-radius:0}.xlHPle .VfPpkd-fmcmS-yrriRe:hover .VfPpkd-fmcmS-OyKIhb::before,.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-fmcmS-OyKIhb::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-fmcmS-OyKIhb::before,.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-fmcmS-OyKIhb::before{transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.xlHPle .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-OyKIhb::before,.xlHPle .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-OyKIhb::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(25,103,210)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(60,64,67)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me){background-color:rgb(241,243,244)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(32,33,36)}.xlHPle .VfPpkd-fmcmS-yrriRe:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(32,33,36)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(25,103,210)}@media all{.GmFilledAutocomplete .mdc-text-field:not(.mdc-text-field--disabled) .mdc-text-field__input::-moz-placeholder{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(95,99,104)}}@media all{.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(95,99,104)}}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(95,99,104)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(60,64,67,.38)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me{background-color:rgba(95,99,104,.04)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(95,99,104,.38)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(95,99,104,.38)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(60,64,67,.38)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgba(95,99,104,.38)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(60,64,67,.38)}@media all{.GmFilledAutocomplete .mdc-text-field.mdc-text-field--disabled .mdc-text-field__input::-moz-placeholder{color:rgba(60,64,67,.38)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(60,64,67,.38)}}@media all{.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(60,64,67,.38)}}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(60,64,67,.38)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(25,103,210)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(197,34,31)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(197,34,31)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(217,48,37)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(197,34,31)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(197,34,31)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(165,14,14)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(165,14,14)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(165,14,14)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(165,14,14)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(25,103,210)}.xlHPle .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(197,34,31)}.xlHPle .VfPpkd-xl07Ob-XxIAqe{box-shadow:0 2px 1px -1px rgba(0,0,0,.2),0 1px 1px 0 rgba(0,0,0,.14),0 1px 3px 0 rgba(0,0,0,.12)}.xlHPle .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:#000;color:var(--mdc-theme-on-surface,#000);position:relative}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(95,99,104)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(60,64,67)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#000;color:var(--mdc-theme-on-surface,#000)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#000;color:var(--mdc-theme-on-surface,#000)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.xlHPle .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}.pxGRyb{display:-moz-inline-box;display:inline-flex;position:relative}.pxGRyb[hidden]{display:none}.pxGRyb .UMrnmb-lP5Lpb-yrriRe,.pxGRyb .UMrnmb-fdMfRe{width:inherit}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px}[dir=rtl] .pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.pxGRyb .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:8px}[dir=rtl] .pxGRyb .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc,.pxGRyb .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:8px;margin-right:0}.pxGRyb .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:48px;padding-right:16px}[dir=rtl] .pxGRyb .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b,.pxGRyb .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:48px}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(60,64,67);color:var(--gm-outlinedtextfield-ink-color,rgb(60,64,67))}.pxGRyb .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(26,115,232);caret-color:var(--gm-outlinedtextfield-caret-color,rgb(26,115,232))}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-helper-text-color,rgb(95,99,104))}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(95,99,104)}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-label-color,rgb(95,99,104))}.pxGRyb .VfPpkd-fmcmS-yrriRe:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(32,33,36)}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(128,134,139);border-color:var(--gm-outlinedtextfield-outline-color,rgb(128,134,139))}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(32,33,36)}@media all{.GmOutlinedAutocomplete .mdc-text-field:not(.mdc-text-field--disabled) .mdc-text-field__input::-moz-placeholder{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-placeholder-color,rgb(95,99,104))}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-placeholder-color,rgb(95,99,104))}}@media all{.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-placeholder-color,rgb(95,99,104))}}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-prefix-color,rgb(95,99,104))}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(95,99,104);color:var(--gm-outlinedtextfield-suffix-color,rgb(95,99,104))}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(95,99,104)}.pxGRyb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(95,99,104)}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-ink-color--disabled,rgba(95,99,104,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(60,64,67,.12);border-color:var(--gm-outlinedtextfield-outline-color--disabled,rgba(60,64,67,.12))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-label-color--disabled,rgba(95,99,104,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(95,99,104,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(95,99,104,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-helper-text-color--disabled,rgba(95,99,104,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-character-counter-color--disabled,rgba(95,99,104,.38))}@media all{.GmOutlinedAutocomplete .mdc-text-field.mdc-text-field--disabled .mdc-text-field__input::-moz-placeholder{color:rgba(60,64,67,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(60,64,67,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(60,64,67,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(60,64,67,.38))}}@media all{.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(60,64,67,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(60,64,67,.38))}}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-prefix-color--disabled,rgba(95,99,104,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(95,99,104,.38);color:var(--gm-outlinedtextfield-suffix-color--disabled,rgba(95,99,104,.38))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(26,115,232);border-color:var(--gm-outlinedtextfield-outline-color--stateful,rgb(26,115,232))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(26,115,232);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(26,115,232))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(217,48,37);caret-color:var(--gm-outlinedtextfield-caret-color--error,rgb(217,48,37))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(217,48,37);color:var(--gm-outlinedtextfield-helper-text-color--error,rgb(217,48,37))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(165,14,14)}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(165,14,14)}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(165,14,14)}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(165,14,14)}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(217,48,37);border-color:var(--gm-outlinedtextfield-outline-color--error,rgb(217,48,37))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(217,48,37);color:var(--gm-outlinedtextfield-icon-color--error,rgb(217,48,37))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(217,48,37);border-color:var(--gm-outlinedtextfield-outline-color--error-stateful,rgb(217,48,37))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(26,115,232);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(26,115,232))}.pxGRyb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(217,48,37);color:var(--gm-outlinedtextfield-label-color--error,rgb(217,48,37))}.pxGRyb .VfPpkd-xl07Ob-XxIAqe{box-shadow:0 2px 1px -1px rgba(0,0,0,.2),0 1px 1px 0 rgba(0,0,0,.14),0 1px 3px 0 rgba(0,0,0,.12);margin-bottom:8px}.pxGRyb.UMrnmb-h0T7hb-OWXEXe-di8rgd-V67aGc .VfPpkd-xl07Ob-XxIAqe,.pxGRyb .VfPpkd-xl07Ob-XxIAqe-OWXEXe-uxVfW-FNFY6c-uFfGwd{margin-bottom:0}.pxGRyb .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:#000;color:var(--mdc-theme-on-surface,#000);position:relative}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(95,99,104)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(60,64,67)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#000;color:var(--mdc-theme-on-surface,#000)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#000;color:var(--mdc-theme-on-surface,#000)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition:opacity .15s linear}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.pxGRyb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}.xQEJ4d .kCI6s{height:3rem}.xQEJ4d .kCI6s .VfPpkd-fmcmS-wGMbrd{font-family:Roboto,Helvetica,Arial,sans-serif;font-size:.875rem}.wlE08e{margin-right:-.25rem}.xQEJ4d .i2Zkcd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me){background-color:rgb(248,249,250)}.xQEJ4d .i2Zkcd.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me{background-color:rgb(248,249,250)}.xQEJ4d .i2Zkcd:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:transparent}.xQEJ4d .i2Zkcd.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:transparent}.xQEJ4d{display:-moz-box;display:flex;position:relative}.xQEJ4d .RSOxzc .VfPpkd-StrnGf-rymPhb{font:.875rem "Roboto",Helvetica,Arial,sans-serif}@keyframes primary-indeterminate-translate{0%{transform:translateX(-145.166611%)}20%{animation-timing-function:cubic-bezier(0.5,0,0.701732,0.495819);transform:translateX(-145.166611%)}59.15%{animation-timing-function:cubic-bezier(0.302435,0.381352,0.55,0.956352);transform:translateX(-61.495191%)}to{transform:translateX(55.444446%)}}@keyframes primary-indeterminate-translate-reverse{0%{transform:translateX(145.166611%)}20%{animation-timing-function:cubic-bezier(0.5,0,0.701732,0.495819);transform:translateX(145.166611%)}59.15%{animation-timing-function:cubic-bezier(0.302435,0.381352,0.55,0.956352);transform:translateX(61.495191%)}to{transform:translateX(-55.4444461%)}}@keyframes primary-indeterminate-scale{0%{transform:scaleX(0.08)}36.65%{animation-timing-function:cubic-bezier(0.334731,0.12482,0.785844,1);transform:scaleX(0.08)}69.15%{animation-timing-function:cubic-bezier(0.06,0.11,0.6,1);transform:scaleX(0.661479)}to{transform:scaleX(0.08)}}@keyframes auxiliary-indeterminate-translate{0%{animation-timing-function:cubic-bezier(0.15,0,0.515058,0.409685);transform:translateX(-54.888891%)}25%{animation-timing-function:cubic-bezier(0.31033,0.284058,0.8,0.733712);transform:translateX(-17.236978%)}48.35%{animation-timing-function:cubic-bezier(0.4,0.627035,0.6,0.902026);transform:translateX(29.497274%)}to{transform:translateX(105.388891%)}}@keyframes auxiliary-indeterminate-translate-reverse{0%{animation-timing-function:cubic-bezier(0.15,0,0.515058,0.409685);transform:translateX(54.888891%)}25%{animation-timing-function:cubic-bezier(0.31033,0.284058,0.8,0.733712);transform:translateX(17.236978%)}48.35%{animation-timing-function:cubic-bezier(0.4,0.627035,0.6,0.902026);transform:translateX(-29.497274%)}to{transform:translateX(-105.388891%)}}@keyframes auxiliary-indeterminate-scale{0%{animation-timing-function:cubic-bezier(0.205028,0.057051,0.57661,0.453971);transform:scaleX(0.08)}19.15%{animation-timing-function:cubic-bezier(0.152313,0.196432,0.648374,1.004315);transform:scaleX(0.457104)}44.15%{animation-timing-function:cubic-bezier(0.257759,0.003163,0.211762,1.38179);transform:scaleX(0.72796)}to{transform:scaleX(0.08)}}@keyframes buffering{to{transform:translateX(-10px)}}@keyframes buffering-reverse{to{transform:translateX(10px)}}@keyframes indeterminate-translate-ie{0%{transform:translateX(-100%)}to{transform:translateX(100%)}}@keyframes indeterminate-translate-reverse-ie{0%{transform:translateX(100%)}to{transform:translateX(-100%)}}.sZwd7c{height:4px;overflow:hidden;position:relative;transform:translateZ(0);transition:opacity 250ms linear;width:100%}.w2zcLc{position:absolute}.xcNBHc,.MyvhI,.l3q5xe{height:100%;position:absolute;width:100%}.w2zcLc{transform-origin:top left;transition:-webkit-transform 250ms ease;transition:transform 250ms ease;transition:transform 250ms ease,-webkit-transform 250ms ease}.MyvhI{transform-origin:top left;transition:-webkit-transform 250ms ease;transition:transform 250ms ease;transition:transform 250ms ease,-webkit-transform 250ms ease;animation:none}.l3q5xe{animation:none}.w2zcLc{background-color:#e6e6e6;height:100%;transform-origin:top left;transition:-webkit-transform 250ms ease;transition:transform 250ms ease;transition:transform 250ms ease,-webkit-transform 250ms ease;width:100%}.TKVRUb{transform:scaleX(0)}.sUoeld{visibility:hidden}.l3q5xe{background-color:#000;display:inline-block}.xcNBHc{background-size:10px 4px;background-repeat:repeat-x;background-image:url('data:image/svg+xml;charset=UTF-8,%3Csvg%20version%3D%271.1%27%20xmlns%3D%27http%3A%2F%2Fwww.w3.org%2F2000%2Fsvg%27%20xmlns%3Axlink%3D%27http%3A%2F%2Fwww.w3.org%2F1999%2Fxlink%27%20x%3D%270px%27%20y%3D%270px%27%20enable-background%3D%27new%200%200%205%202%27%20xml%3Aspace%3D%27preserve%27%20viewBox%3D%270%200%205%202%27%20preserveAspectRatio%3D%27none%20slice%27%3E%3Ccircle%20cx%3D%271%27%20cy%3D%271%27%20r%3D%271%27%20fill%3D%27%23e6e6e6%27%2F%3E%3C%2Fsvg%3E');visibility:hidden}.sZwd7c.B6Vhqe .MyvhI{transition:none}.sZwd7c.B6Vhqe .TKVRUb{animation:primary-indeterminate-translate 2s infinite linear}.sZwd7c.B6Vhqe .TKVRUb>.l3q5xe{animation:primary-indeterminate-scale 2s infinite linear}.sZwd7c.B6Vhqe .sUoeld{animation:auxiliary-indeterminate-translate 2s infinite linear;visibility:visible}.sZwd7c.B6Vhqe .sUoeld>.l3q5xe{animation:auxiliary-indeterminate-scale 2s infinite linear}.sZwd7c.B6Vhqe.ieri7c .l3q5xe{transform:scaleX(0.45)}.sZwd7c.B6Vhqe.ieri7c .sUoeld{animation:none;visibility:hidden}.sZwd7c.B6Vhqe.ieri7c .TKVRUb{animation:indeterminate-translate-ie 2s infinite ease-out}.sZwd7c.B6Vhqe.ieri7c .TKVRUb>.l3q5xe,.sZwd7c.B6Vhqe.ieri7c .sUoeld>.l3q5xe{animation:none}.sZwd7c.juhVM .w2zcLc,.sZwd7c.juhVM .MyvhI{right:0;transform-origin:center right}.sZwd7c.juhVM .TKVRUb{animation-name:primary-indeterminate-translate-reverse}.sZwd7c.juhVM .sUoeld{animation-name:auxiliary-indeterminate-translate-reverse}.sZwd7c.juhVM.ieri7c .TKVRUb{animation-name:indeterminate-translate-reverse-ie}.sZwd7c.qdulke{opacity:0}.sZwd7c.jK7moc .sUoeld,.sZwd7c.jK7moc .TKVRUb,.sZwd7c.jK7moc .sUoeld>.l3q5xe,.sZwd7c.jK7moc .TKVRUb>.l3q5xe{animation-play-state:paused}.sZwd7c.D6TUi .xcNBHc{animation:buffering 250ms infinite linear;visibility:visible}.sZwd7c.D6TUi.juhVM .xcNBHc{animation:buffering-reverse 250ms infinite linear}.d1dlne,.Ax4B8{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1;-moz-box-flex:1;flex:1}.L6J0Pc{-moz-box-flex:1;-moz-box-flex:1;flex:1}.v5yLH,.v5yLH .d1dlne,.v5yLH .Ax4B8{display:inline}.BBOA1c{position:absolute;height:4px;bottom:1px;left:1px;right:1px;overflow-x:hidden;background-color:#fff;display:none}.L6J0Pc.ge6pde .BBOA1c{display:block}.u3WVdc{position:absolute;right:0;left:0;z-index:1;outline:none;overflow-y:auto}.u3WVdc[data-childcount="0"],.u3WVdc[data-expanded=false]{display:none}.Cigftf{position:relative;top:-24px}.Ax4B8{position:relative}.yNVtPc{position:absolute;left:0;width:100%;opacity:.3}.Ax4B8,.yNVtPc{background-color:transparent;color:inherit;font:inherit;line-height:inherit}.Ax4B8::-ms-clear{display:none}.d1dlne,.Ax4B8,.yNVtPc{height:100%}.umNhxf{overflow-x:hidden;text-overflow:ellipsis;white-space:nowrap}.MkjOTb{cursor:default}.VOEIyf,.VOEIyf .jBmls,.oKubKe{font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;color:#222}.VOEIyf{display:inline-block;height:34px;line-height:34px}.IjMZm{display:inline-block;height:auto;line-height:auto}.VOEIyf .ZAGvjd{border-color:transparent;border-style:solid;border-width:0 1px;outline:none}.oKubKe,.VOEIyf .ZAGvjd{-moz-box-sizing:border-box;box-sizing:border-box;padding:0 16px}.VOEIyf .jBmls{-moz-box-sizing:border-box;box-sizing:border-box;padding:8px 0;border:1px solid rgba(0,0,0,.2);background-color:#fff;-moz-border-radius:0 0 2px 2px;border-radius:0 0 2px 2px;-moz-box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2)}.oKubKe{line-height:40px}.oKubKe[aria-selected=true]{background-color:#eee}.oKubKe.RDPZE{color:rgba(0,0,0,.38)}.SmXtye{margin:7px 0;border-top:1px solid #dadada}.D4D33b{overflow-x:hidden;text-overflow:ellipsis;white-space:nowrap}.uVccjd{box-flex:0;flex-grow:0;-moz-user-select:none;-moz-transition:border-color .2s cubic-bezier(0.4,0,0.2,1);transition:border-color .2s cubic-bezier(0.4,0,0.2,1);border:10px solid rgba(0,0,0,.54);-moz-border-radius:3px;border-radius:3px;-moz-box-sizing:content-box;box-sizing:content-box;cursor:pointer;display:inline-block;max-height:0;max-width:0;outline:none;overflow:visible;position:relative;vertical-align:middle;z-index:0}.uVccjd.ZdhN5b{border-color:rgba(255,255,255,.7)}.uVccjd.ZdhN5b[aria-disabled=true]{border-color:rgba(255,255,255,.3)}.uVccjd[aria-disabled=true]{border-color:#bdbdbd;cursor:default}.uHMk6b{-moz-transition:all .1s .15s cubic-bezier(0.4,0,0.2,1);transition:all .1s .15s cubic-bezier(0.4,0,0.2,1);-moz-transition-property:transform,border-radius;transition-property:transform,border-radius;border:8px solid white;left:-8px;position:absolute;top:-8px}[aria-checked=true]>.uHMk6b,[aria-checked=mixed]>.uHMk6b{-moz-transform:scale(0);transform:scale(0);transition:-webkit-transform .1s cubic-bezier(0.4,0,0.2,1);transition:transform .1s cubic-bezier(0.4,0,0.2,1);transition:transform .1s cubic-bezier(0.4,0,0.2,1),-webkit-transform .1s cubic-bezier(0.4,0,0.2,1);-moz-border-radius:100%;border-radius:100%}.B6Vhqe .TCA6qd{left:5px;top:2px}.N2RpBe .TCA6qd{left:10px;-moz-transform:rotate(-45deg);transform:rotate(-45deg);-moz-transform-origin:0;transform-origin:0;top:7px}.TCA6qd{height:100%;pointer-events:none;position:absolute;width:100%}.rq8Mwb{-moz-animation:quantumWizPaperAnimateCheckMarkOut .2s forwards;animation:quantumWizPaperAnimateCheckMarkOut .2s forwards;clip:rect(0,20px,20px,0);height:20px;left:-10px;position:absolute;top:-10px;width:20px}[aria-checked=true]>.rq8Mwb,[aria-checked=mixed]>.rq8Mwb{-moz-animation:quantumWizPaperAnimateCheckMarkIn .2s .1s forwards;animation:quantumWizPaperAnimateCheckMarkIn .2s .1s forwards;clip:rect(0,20px,20px,20px)}@media print{[aria-checked=true]>.rq8Mwb,[aria-checked=mixed]>.rq8Mwb{clip:auto}}.B6Vhqe .MbUTNc{display:none}.MbUTNc{border:1px solid #fff;height:5px;left:0;position:absolute}.B6Vhqe .Ii6cVc{width:8px;top:7px}.N2RpBe .Ii6cVc{width:11px}.Ii6cVc{border:1px solid #fff;left:0;position:absolute;top:5px}.PkgjBf{-moz-transform:scale(2.5);transform:scale(2.5);-moz-transition:opacity 0.15s ease;transition:opacity 0.15s ease;background-color:rgba(0,0,0,0.2);-moz-border-radius:100%;border-radius:100%;height:20px;left:-10px;opacity:0;outline:.1px solid transparent;pointer-events:none;position:absolute;top:-10px;width:20px;z-index:-1}.ZdhN5b .PkgjBf{background-color:rgba(255,255,255,0.2)}.qs41qe>.PkgjBf{-moz-animation:quantumWizRadialInkSpread .3s;animation:quantumWizRadialInkSpread .3s;animation-fill-mode:forwards;opacity:1}.i9xfbb>.PkgjBf{background-color:rgba(0,150,136,0.2)}.u3bW4e>.PkgjBf{-moz-animation:quantumWizRadialInkFocusPulse .7s infinite alternate;animation:quantumWizRadialInkFocusPulse .7s infinite alternate;background-color:rgba(0,150,136,0.2);opacity:1}@keyframes quantumWizPaperAnimateCheckMarkIn{0%{clip:rect(0,0,20px,0)}to{clip:rect(0,20px,20px,0)}}@keyframes quantumWizPaperAnimateCheckMarkOut{0%{clip:rect(0,20px,20px,0)}to{clip:rect(0,20px,20px,20px)}}.aiSeRd{border-color:#5f6368}.aiSeRd:before{bottom:-24px;content:"";display:block;height:48px;left:-24px;position:absolute;right:-24px;top:-24px;width:48px}.aiSeRd.N2RpBe,.aiSeRd.B6Vhqe{border-color:#1a73e8}.aiSeRd.RDPZE{border-color:#bdc1c6}.aiSeRd>.MbhUzd{height:16px;width:16px;left:-8px;top:-8px}.aiSeRd:hover>.MbhUzd{-moz-animation:quantumWizRadialInkSpread;animation:quantumWizRadialInkSpread;animation-fill-mode:forwards;background-color:rgba(32,33,36,0.039)}.aiSeRd.N2RpBe:hover>.MbhUzd{background-color:rgba(26,115,232,0.039)}.aiSeRd:focus>.MbhUzd{-moz-animation:quantumWizRadialInkSpread;animation:quantumWizRadialInkSpread;animation-fill-mode:forwards;background-color:rgba(32,33,36,0.078)}.aiSeRd.N2RpBe:focus>.MbhUzd{background-color:rgba(26,115,232,0.078)}.aiSeRd.RDPZE:focus>.MbhUzd,.aiSeRd.RDPZE:hover>.MbhUzd{display:none}.aiSeRd.u3bW4e>.MbhUzd{-moz-animation:quantumWizRadialInkSpread;animation:quantumWizRadialInkSpread;animation-fill-mode:forwards;background-color:rgba(32,33,36,0.122)}.aiSeRd.N2RpBe.u3bW4e>.MbhUzd{background-color:rgba(26,115,232,0.122)}.aiSeRd.qs41qe>.MbhUzd{-moz-animation:quantumWizRadialInkFocusPulse .3s;animation:quantumWizRadialInkFocusPulse .3s;animation-fill-mode:forwards;background-color:rgba(32,33,36,0.161)}.aiSeRd.N2RpBe.qs41qe>.MbhUzd{background-color:rgba(26,115,232,0.161)}.gj14oe:hover>.MbhUzd{-moz-animation:quantumWizRadialInkSpread;animation:quantumWizRadialInkSpread;animation-fill-mode:forwards;background-color:rgba(255,255,255,0.078)}.gj14oe:focus>.MbhUzd{-moz-animation:quantumWizRadialInkSpread;animation:quantumWizRadialInkSpread;animation-fill-mode:forwards;background-color:rgba(255,255,255,0.161)}.gj14oe.RDPZE:hover>.MbhUzd{display:none}.gj14oe.u3bW4e>.MbhUzd{-moz-animation:quantumWizRadialInkSpread;animation:quantumWizRadialInkSpread;animation-fill-mode:forwards;background-color:rgba(255,255,255,0.239)}.gj14oe.qs41qe>.MbhUzd{-moz-animation:quantumWizRadialInkFocusPulse .3s;animation:quantumWizRadialInkFocusPulse .3s;animation-fill-mode:forwards;background-color:rgba(255,255,255,0.322)}.BIHLNc{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.aiSeRd+.Mk3P9d{margin-left:8px}.aiSeRd.RDPZE+.Mk3P9d{color:rgba(0,0,0,.38)}.mSdN4b{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-flow:column wrap;max-width:100%}@charset "UTF-8";.odb4eb{border-bottom:.0625rem solid;color:rgb(218,220,224);margin-bottom:.5rem}.qiFkmc .VfPpkd-TkwUic{height:52px;display:-moz-box;display:flex;-moz-box-align:baseline;align-items:baseline}.qiFkmc .VfPpkd-TkwUic::before{display:inline-block;width:0;height:40px;content:"";vertical-align:0}.qiFkmc.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS::before{content:"​"}.qiFkmc.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS-haAclf{height:100%;display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center}.qiFkmc.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic::before{display:none}.qiFkmc .VfPpkd-t08AT-Bz112c{width:20px;height:20px}.qiFkmc.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{max-width:calc(100% - 60px)}.qiFkmc.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:calc(133.3333333333% - 80px)}.qiFkmc .VfPpkd-StrnGf-rymPhb-ibnC6b,.qiFkmc .VfPpkd-aJasdd-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:44px}.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:60px}.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-Gtdoyb{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-pack:center;justify-content:center}.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS{margin-top:0;margin-bottom:0;line-height:1.4}.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS::before,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS::after{display:none}.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.qiFkmc .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:68px}.qiFkmc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-TkwUic{background-color:rgb(248,249,250)}.qiFkmc .VfPpkd-OkbHre .VfPpkd-rymPhb-fpDzbe-fmcmS{font-size:14px}.qiFkmc .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-width:0}.qiFkmc .VfPpkd-uusGie-fmcmS{font-size:14px}.Y7l6jd{width:100%}.XxyAsb{background:url('https://www.gstatic.com/docs/doclist/images/mediatype/icon_1_document_x64.png') center no-repeat}.qurv4d{background:url('https://www.gstatic.com/docs/doclist/images/mediatype/icon_1_presentation_x64.png') center no-repeat}.teCq2b{background:url('https://www.gstatic.com/docs/doclist/images/mediatype/icon_1_sheets_x64.png') center no-repeat}.O1YELb{background:url('https://www.gstatic.com/docs/doclist/images/mediatype/icon_1_drawing_x64.png') center no-repeat}.aV9qc{background:url('https://www.gstatic.com/docs/doclist/images/mediatype/icon_2_form_x64.png') center no-repeat}.XxyAsb,.qurv4d,.teCq2b,.O1YELb,.aV9qc{background-size:contain;height:1.25rem;width:1.25rem}.mMfeif.ubvFYc{line-height:2rem;margin-left:1rem}.moEOjf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-shrink:0}.TDK0Zb{align-items:stretch;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;box-flex:1;flex-grow:1}.svNSpd{border-color:#e8eaed;-moz-border-radius:50%;border-radius:50%;border-style:solid;border-width:0.0625rem;height:3rem;margin:0.5rem;margin-bottom:0.5rem;width:3rem}.yKnF7e{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;margin-right:0.0625rem}.rkHJle .Ce1Y1c{opacity:1}.a7AG0{height:1.125rem;width:1.125rem}.zAg7wc{font-size:1.25rem;height:1.25rem;width:1.25rem}.qYr7gb{-moz-column-gap:0.875rem;column-gap:0.875rem;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:wrap;flex-wrap:wrap}.gPDsDb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;margin-top:0.25rem;max-height:13.75rem;overflow:auto;padding-bottom:1rem;padding-right:1.5rem}.i3bmcb{border-color:#e8eaed;-moz-border-radius:50%;border-radius:50%;border-style:solid;border-width:0.0625rem;height:3rem;margin:0.75rem;margin-bottom:0.5rem;width:3rem}.SwCXPc{letter-spacing:.01785714em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;font-weight:500;line-height:1.25rem;margin-bottom:0.875rem;max-width:4.625rem;text-align:center;word-wrap:break-word}.lrj7Bb:focus{border:0.125rem solid #185abc;-moz-border-radius:0.375rem;border-radius:0.375rem}.Tjbfle{letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:.75rem;font-weight:400;-moz-border-radius:3.25rem;border-radius:3.25rem;color:white;line-height:1.25rem;padding:0 0.375rem;position:absolute;right:-1.5rem}.RWzxl{-moz-user-select:none;-moz-user-select:none;display:inline-block;outline:none;width:200px}.KzNPgc{position:relative;vertical-align:top}.JGptt{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.Hvn9fb{-moz-box-flex:1;box-flex:1;flex-grow:1;flex-shrink:1;background-color:transparent;border:none;display:block;font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;margin:0;min-width:0%;outline:none;padding:.125em 0;z-index:0}.SPcBRc{background-color:rgba(0,0,0,.12);height:1px;margin:0;padding:0;width:100%}.kPBwDb{transform:scaleX(0);background-color:#03a9f4;height:2px;margin:0;padding:0;width:100%}.RWzxl.RDPZE .Hvn9fb{color:rgba(0,0,0,.38)}.RWzxl.RDPZE>.KzNPgc>.SPcBRc{background:none;border-bottom:1px dotted rgba(0,0,0,.38)}.kPBwDb.Y2Zypf{animation:quantumWizSimpleInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1)}.RWzxl.u3bW4e>.KzNPgc>.kPBwDb{animation:quantumWizSimpleInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);transform:scaleX(1)}.BYyR7e{color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;max-width:100%;overflow:hidden;pointer-events:none;position:absolute;text-overflow:ellipsis;white-space:nowrap}.RWzxl.CDELXb>.KzNPgc>.BYyR7e{display:none}@keyframes quantumWizSimpleInputRemoveUnderline{0%{transform:scaleX(1);opacity:1}to{transform:scaleX(1);opacity:0}}@keyframes quantumWizSimpleInputAddUnderline{0%{transform:scaleX(0)}to{transform:scaleX(1)}}.V6WXSe{-moz-box-align:center;box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;font-size:13px;font-weight:400;min-height:48px}.V6WXSe .mIZh1c{margin-top:4px;visibility:hidden}.V6WXSe:hover .mIZh1c,.W0RsD.u3bW4e .mIZh1c{visibility:visible}.EsoU5c{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-align:center;box-align:center;align-items:center;flex-shrink:0}.UhHij{margin-right:12px}.QxM9Wc{opacity:.5}.NreIxc{width:48px}.W0RsD{width:100%}.W0RsD input{font-size:13px;width:100%}.uEtsdd{margin-top:8px;min-width:0;box-flex:1;flex-grow:1}.uEtsdd.xkhr8{box-flex:0;flex-grow:0;margin-right:4px}.uEtsdd.xkhr8 .snByac{color:rgba(0,0,0,.54);font-size:13px;position:static}.xkhr8 input{cursor:pointer;position:absolute;top:0}.cy9MSc{color:#4285f4;cursor:pointer;font-weight:500;margin-left:4px;text-align:center;text-transform:uppercase}.yrhGr{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-align:center;box-align:center;align-items:center;box-flex:1;flex-grow:1}.si40te{height:24px;visibility:hidden;width:42px}.V6WXSe:hover .si40te{visibility:visible}.CCJ0ld-Jup3Tc .si40te,.dgl2Hf .V6WXSe.IwUXg .si40te{visibility:visible}.CCJ0ld-Jup3Tc .yrhGr{-moz-box-shadow:0px 1px 1px 0px rgba(0,0,0,.14),0px 2px 1px -1px rgba(0,0,0,.12),0px 1px 3px 0px rgba(0,0,0,.2);box-shadow:0px 1px 1px 0px rgba(0,0,0,.14),0px 2px 1px -1px rgba(0,0,0,.12),0px 1px 3px 0px rgba(0,0,0,.2);background:#fff;opacity:.7}.si40te .QNGjdb-zJVW9d{cursor:move;text-align:center;opacity:.3}.Kq74Wb{margin:-0.5rem -1rem 0;padding-bottom:1rem;overflow:hidden}.Kq74Wb .W0RsD input,.Kq74Wb .xkhr8 .snByac{font-size:0.875rem}.OA0qNb .bpT8Rd{display:none}.GtIyje{color:#b31412}.RdbXWd{height:0.625rem}.j1BhHb{line-height:1;padding:0.5rem 0}.kCyxtd.RDPZE .j1BhHb{color:rgba(68,68,68,0.502);cursor:default}.JPdR6b.e5Emjc .nwYmvb.z80M1{padding-left:3.5rem;padding-right:1rem}.nwYmvb{flex-flow:column nowrap}.nwYmvb .PCdOIb{height:100%;left:1rem}.nwYmvb .uyYuVb{font-size:0.8125rem;height:auto;line-height:1.25rem}.FAVvUd.z80M1.N2RpBe:before{content:none}.FAVvUd .nIu6nb{background-position:-13.25rem 0;height:1.5rem;width:1.5rem}.FAVvUd.N2RpBe .nIu6nb{background-position:-13.25rem -2.5rem;height:1.5rem;width:1.5rem}.wbGyrc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-flow:column;height:3.5rem;justify-content:center;width:7.5rem}.kuntz{flex-shrink:0;margin-right:1rem}.apMwAf{text-overflow:ellipsis;overflow:hidden;white-space:nowrap}.bUqWxf{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;color:rgba(0,0,0,.549)}.EKkFUc .wbGyrc{color:rgba(0,0,0,.549)}.EKkFUc .bUqWxf{color:rgba(0,0,0,.38)}@media (max-width:40em){.oCUiN .j1BhHb,.nwYmvb .uyYuVb{font-size:0.875rem}}.HMUCnd{width:100%}.xe721c{color:rgba(0,0,0,.549)}.HMUCnd .LMgvRb .oJeWuf,.HMUCnd .OA0qNb .oJeWuf{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;display:block}.J1NSgc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row}.QTi9Ve{padding:0.0625rem;margin-left:0.5rem;margin-right:0.5rem;height:fit-content;align-self:center;margin-bottom:0.5rem}@media (max-width:40em){.HMUCnd .LMgvRb .oJeWuf{font-size:0.875rem}}.zYkTW{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.GV4Keb{height:3rem;margin-bottom:0;margin-top:0;width:100%}.JbvUD{max-height:31.25rem}.DHnzaf{visibility:hidden}.RDGyy{height:3rem;width:100%}.qbzgQb{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-pack:justify;justify-content:space-between;margin-bottom:.75rem}.uHsvzf{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:500}.KDyM1e{margin-left:1.75rem;max-width:14.25rem}.O98Lj{color:#333;font-family:"Roboto",Helvetica,Arial,sans-serif;font-size:0.8125rem;line-height:1.25rem;position:relative}.QTMzUe{border:none;outline:none;width:100%}input.QTMzUe::-webkit-input-placeholder,input.QTMzUe:-moz-placeholder,input.QTMzUe::-moz-placeholder,input.QTMzUe:-ms-input-placeholder{color:rgba(0,0,0,.24)}input.QTMzUe:disabled{background-color:#f5f5f5}.Yiql6e p{margin:0}.Lzdwhd-BrZSOd{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;-moz-user-select:none;color:rgba(0,0,0,.24);position:absolute}.Lzdwhd-AyKMt{border-bottom:0.0625rem solid rgba(0,0,0,.24);padding-bottom:0.0625rem}.Lzdwhd-AyKMt:focus{border-bottom:#377dfa solid 0.125rem;padding-bottom:0}.QTMzUe{box-sizing:border-box;padding:0.875rem}.QTMzUe:focus{border-bottom-width:0.125rem;border-bottom-style:solid;padding-bottom:0.75rem}.Lzdwhd-AyKMt.iTy5c{border:none}.Lzdwhd-AyKMt{cursor:text;outline:none;position:relative;word-wrap:break-word;min-height:1.25rem}@media (max-width:40em){.O98Lj{font-size:0.875rem}}.ztA2jd-auswjd{background-color:#eee}.ztA2jd-SUR3Rd{-moz-box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);box-shadow:0 0.0625rem 0.125rem rgba(0,0,0,.12),0 0 0.0625rem rgba(0,0,0,.12);background:#fff;box-sizing:border-box;font-family:"Roboto",Helvetica,Arial,sans-serif;font-size:0.8125rem;position:absolute;z-index:1192}.ztA2jd-oKdM2c{box-sizing:border-box;line-height:1.75rem;height:3rem;padding:0.5rem 1rem;width:100%}.f68nG{font-weight:500}.aIx74 .snByac{white-space:nowrap}.aIx74 .DPvwYc{display:inline-block;color:#9e9e9e;pointer-events:none;vertical-align:middle;margin:-0.25rem 0}.aIx74 .RDPZE .DPvwYc{color:#bdbdbd}.olCKnc{flex-shrink:0}.BUagKb{display:inline-block;min-width:2.5rem;text-transform:none}.RDPZE .BUagKb{color:inherit}.y2d25{background-color:#fff;-moz-box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);box-shadow:0px 8px 10px 1px rgba(0,0,0,.14),0px 3px 14px 2px rgba(0,0,0,.12),0px 5px 5px -3px rgba(0,0,0,.2);-moz-border-radius:4px;border-radius:4px;position:absolute;width:16.25rem;z-index:1200}.ECK80e{border-bottom:0.0625rem solid #e0e0e0;cursor:default;font-size:0.9375rem;padding:1rem 1.5rem}.DTnYMd{padding:1.5rem}.gA55mc{margin-bottom:1rem}@media (max-width:40em){.aIx74{font-size:0.875rem}.ECK80e{font-size:1rem}}.dKKcxf,.STMvPe{background:#f8f9fa;cursor:pointer;margin-bottom:0.5rem}input.tAUuQ{background:transparent}input.tAUuQ:disabled{background:transparent;color:rgba(0,0,0,.549)}input.tAUuQ:disabled+.XOaaUb{color:#bdbdbd}.RPt7lf{position:relative}.dKKcxf input.tAUuQ:not(:disabled){cursor:pointer}.STMvPe{margin-top:1rem}.XOaaUb{pointer-events:none}.Y6kebb,.XOaaUb{cursor:pointer;opacity:0.54;position:absolute}.Y6kebb,.XOaaUb{right:0.875rem;top:0.75rem}.Y6kebb{color:#5f6368}.NE9bBb{background:#f8f9fa;box-sizing:border-box;color:rgba(0,0,0,.549)!important;padding:0.875rem;width:100%}.NE9bBb:focus,.a2YH8d .NE9bBb,.a2YH8d input.tAUuQ{border-bottom:0.125rem solid rgba(0,0,0,.24);padding-bottom:0.75rem}.a2YH8d .NE9bBb,.a2YH8d .NE9bBb:focus,.a2YH8d input.tAUuQ{border-color:#ea4335!important}.SQJ88{color:#ea4335;font-size:0.75rem;margin-top:0.25rem}.aK5JE .RPt7lf,.fEejq:not(.a2YH8d) .SQJ88,.RPt7lf:not(.miHM0e)>.tAUuQ,.RPt7lf:not(.miHM0e) .Y6kebb,.RPt7lf.miHM0e>.NE9bBb,.RPt7lf.miHM0e:not(.Y5OfKb)>.XOaaUb,.RPt7lf.dKKcxf:not(.miHM0e)+.RPt7lf.STMvPe{display:none}@media (max-width:40em){.fEejq,.tAUuQ{font-size:0.875rem}}.Rt2Mob{height:3rem;padding:0 1.5rem}.SQM07d,.IfzqGf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;width:100%}.TIKlJe .hqBSCb .VfPpkd-TkwUic{background-color:#f8f9fa;height:3rem}.TIKlJe{width:100%}.TIKlJe .LMgvRb .oJeWuf,.TIKlJe .OA0qNb .oJeWuf{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;display:block}.a4Vkrf{min-width:15rem}.c8GN4d{max-height:18.75rem}@media (max-width:40em){.TIKlJe .LMgvRb .oJeWuf{font-size:0.875rem}.a4Vkrf{min-width:25rem}}.sRTzRd .oJeWuf{height:3rem}.sRTzRd .mIZh1c{display:none}.wc5HEf{height:1.5rem;opacity:0.54;width:1.5rem}.bDkUbc{border-bottom-style:solid;border-bottom-width:0.0625rem;color:#dadce0}.AysVpb .VfPpkd-OkbHre .VfPpkd-rymPhb-fpDzbe-fmcmS{font-size:14px}.AysVpb .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-width:0}.AysVpb .VfPpkd-uusGie-fmcmS{font-size:14px}.h4f0L{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row}.pe3QUd{-moz-box-flex:1;flex-grow:1}.Isz4Oc{color:rgb(95,99,104)}.nNvQ{color:rgb(154,160,166)}.KEwy9{text-overflow:ellipsis;overflow:hidden;white-space:nowrap}.pvb7Pc{border-bottom:0.0625rem solid #e0e0e0;height:3.5rem;padding-right:0.5rem;white-space:nowrap}.YXgoed{color:#fff;cursor:default;flex-shrink:0;height:3.5rem;line-height:0;width:3.5rem}.hgjBDc{background-color:#fff;overflow:hidden;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.hgjBDc .YioO4d{margin-bottom:0}.LZqXdf{-moz-box-flex:1 1 auto;flex:1 1 auto;padding-top:1.5rem;overflow-y:auto}.aqlftc{margin:0 1.5rem 1.5rem}.AWfQId{-moz-flex-wrap:wrap;flex-wrap:wrap;padding:0 0.5rem 0.5rem 1.5rem}.AWfQId>*,.rxO3db>*{flex-shrink:0}.w1v75b{box-flex:99999;flex-grow:99999}.AWfQId .w1v75b,.AWfQId .rxO3db{margin-bottom:1rem;margin-right:1rem}.AWfQId .QqqDDf{height:3rem}.rxO3db{box-flex:1;flex-grow:1;justify-content:flex-end}@media (max-width:30em){.AWfQId .w1v75b{-moz-flex-wrap:wrap;flex-wrap:wrap;max-width:18.75rem}}.TQX6ub:not(:empty){margin-bottom:1.5rem;padding:0 1.5rem}.KbjbQd{-moz-box-flex:0 0 auto;flex:0 0 auto}@media (max-width:40em){.TQX6ub:not(:empty){margin-bottom:1rem}}.p9YKmd.p9YKmd{margin-right:0.5rem}.mpfp4{margin-right:1.5rem}@media not all and (max-width:40em){.tS2rsb{display:none}.IL2Cre{align-items:stretch;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;box-flex:1;flex-grow:1;margin:-1rem 0.5rem}.hja3X{border-right:0.0625rem solid #e0e0e0;box-flex:1;flex-grow:1;min-width:0;padding:1.5rem;padding-left:0;padding-bottom:0.5rem}.TdC1bb{background-color:#f8f9fa;margin-left:-1.5rem;padding-left:1.5rem}.NVmm2e{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center}.Sl8ssb{box-sizing:border-box;margin-bottom:1.5rem;min-width:0;overflow:visible;padding:1.5rem;padding-bottom:0.5rem;width:60rem}.uWetjb{flex-shrink:0;padding:1.5rem 0;padding-left:1.5rem}}@media (max-width:40em){.Sl8ssb{margin-bottom:1.5rem;overflow:visible;padding:1.25rem 0.875rem 0.875rem 0.875rem}.uWetjb{margin-bottom:2.5rem}.IY1wn{display:none}}@media not all and (max-width:900px){.XZDC9d{max-width:60rem;align-items:stretch;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;box-flex:1;flex-grow:1;margin-bottom:1.5rem}.bGJJfc{border-right:0.0625rem solid #e0e0e0}}@media (max-width:900px){.XZDC9d{box-flex:1;flex-grow:1;margin-bottom:1.5rem}.bGJJfc{border-bottom:0.0625rem solid #e0e0e0}}.ThlZVb{box-flex:1;flex-grow:1;padding-top:1rem;padding-left:1.5rem}.Ocq0Sc{box-sizing:border-box;box-flex:0;flex-grow:0;min-width:14.375rem}.AUczsd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.PyxdTe{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:1;flex-grow:1;padding:0.875rem 1.5rem}.X6EBqc,.QwKx3b{align-items:center;color:#5f6368;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;margin-right:0.25rem}.tzhXFf{margin:-0.75rem 0.5rem 0}@media (min-width:1152px){.Ocq0Sc{width:20.625rem}}.AOhYp{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-bottom:1rem;overflow:hidden}.qASq1{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:1;flex-grow:1;-moz-flex-wrap:wrap;flex-wrap:wrap}.AOhYp .AHfDQd{box-flex:1;flex-grow:1;min-width:0}.TWyWEc{margin-left:1rem}.czCkDc{border-top:0.0625rem solid #e0e0e0;margin:0 -1rem 1.5rem}.Qupzef{margin-bottom:1rem}@media not all and (max-width:40em){.AJRyDb{margin-left:3rem}}@media (max-width:900px){.jVw62e{width:100%}.TWyWEc{box-flex:1;flex-grow:1;margin-left:0;margin-top:1rem}}.ec5iTb{margin:-1.5rem;margin-bottom:1.5rem}@media (max-width:40em){.ec5iTb{margin:-1rem -1rem 1.5rem}}.YioO4d{margin-bottom:1rem;width:9.375rem}.uWetjb .LMgvRb{min-width:0}@media (min-width:780px){.YioO4d.hioilb{width:19.75rem}}@media (max-width:40em),(min-width:780px){.CWm61{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.CWm61 .YioO4d+.YioO4d{margin-left:1rem}}.u8xvqb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.u8xvqb .YioO4d+.YioO4d{margin-left:1rem}@media (max-width:40em){.YioO4d{width:-moz-calc((100% - 1rem)/2);width:calc((100% - 1rem)/2)}.YioO4d.hioilb{width:100%}}.gtuckc{margin-bottom:0.5rem}.X4Eo2e{width:44px;height:44px;padding:11px;font-size:22px}.X4Eo2e svg,.X4Eo2e img{width:22px;height:22px}.xS05rc{width:44px;height:44px;padding:11px;font-size:22px}.xS05rc svg,.xS05rc img{width:22px;height:22px}.vmQOqd{color:rgb(232,234,237);margin-bottom:.75rem}.NaHd8c{margin-left:-.9375rem;margin-bottom:-.9375rem}.CWm61{-moz-box-align:end;align-items:flex-end}.S51BW .KRoqRc{min-height:6.25rem}.w1NASc{padding:.3125rem 0;width:100%}.w1NASc .eU809d{top:1.625rem}.w1NASc .LMgvRb{max-width:100%}.cZSNUb{margin-bottom:0.5rem}.MGjN3e{min-height:2.125rem}.MGjN3e .LsSwGf{margin-right:0.5rem}.ZZAGKd .bEd2J{margin-bottom:.875rem;margin-top:.875rem}.zOtZye{min-height:4.5rem}.zTrXGf{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:100%;position:relative;z-index:0}.qk0lee{cursor:pointer;box-flex:1;flex-grow:1}.qk0lee:focus:after{background:#f5f5f5;content:"";height:100%;left:0;position:absolute;top:0;width:100%;z-index:-1}.qk0lee:hover .K6Ovqd{color:inherit}.U2zcIf{margin-left:0.5rem;padding:1rem}.fidHdf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-left:1rem;padding:0 0.75rem}.K6Ovqd{align-items:center;color:rgba(0,0,0,.549);display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1 1 auto;flex:1 1 auto;height:100%;justify-content:flex-start}.Bw8p0d .KbjbQd{display:none;padding-top:1.5rem}.H87RP{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;margin-top:4rem;text-align:center}.H87RP img{margin-bottom:1.5rem;max-width:25vw}.CMXcoc{padding:1.5rem}.CMXcoc .z3vRcc{margin-bottom:.5rem}.y9k09d:not(:empty){margin-top:1.5rem}.MdjMac{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;padding:2rem 1rem 2rem 2rem}@media (max-width:30rem){.MdjMac{-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;padding:2rem 1rem;text-align:center}}.Fnu4gf{flex-shrink:0;height:5.625rem;margin-right:2.5rem}@media (max-width:30rem){.Fnu4gf{margin-bottom:1rem}}.B14Gwb{display:-moz-box;display:flex;-moz-box-pack:end;justify-content:end;margin-top:.5rem}@media (max-width:30rem){.B14Gwb{display:block;margin-top:1rem}}.aQkHxe{margin-bottom:.5rem}.kDu3nf{height:9.375rem;margin-top:4rem}.n86u6b{margin:2.1875rem 0 1rem 0;width:16.625rem}.erXmAf{margin-right:1rem}.xPAMbf{align-items:center;border-bottom:0.0625rem solid #e0e0e0;box-sizing:border-box;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;height:3.75rem;padding:0.5rem 1.5rem 0.5rem 1.5rem;position:relative}.UvQypf.xPAMbf{cursor:pointer}.WaqnWd{align-items:center;box-sizing:border-box;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:0 0 auto;flex:0 0 auto;height:2.25rem;justify-content:center;margin-right:1rem;width:2.25rem}.cQaDA{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1 1 auto;flex:1 1 auto;flex-direction:row;overflow:hidden}.ToDHyd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1 1 auto;flex:1 1 auto;flex-direction:row;overflow:hidden;flex-direction:column}.Wd54if{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:0 0 auto;flex:0 0 auto}.k19Ou,.Jd0Ule{box-sizing:border-box;-moz-box-flex:0 0 auto;flex:0 0 auto;margin-left:0.5rem;margin-right:-1rem;width:2.5rem}.xPAMbf .ptXozb{bottom:0;left:0;position:absolute;right:0;top:0;z-index:-1}.SPoV1e{box-sizing:border-box;padding:1rem 1.5rem 1rem 1.5rem;width:100%}.tmJXcf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.aKNfrc{margin-top:1rem;margin-bottom:-0.5rem}.yJz7Ve{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1 1 auto;flex:1 1 auto;flex-direction:column;overflow:hidden}.HfeSwf{-moz-box-flex:0 0 auto;flex:0 0 auto;margin-left:1rem}.stPFhf{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;justify-content:space-between}@media (max-width:40em){.tmJXcf{flex-direction:column}.yJz7Ve+.HfeSwf{margin-top:1rem}.HfeSwf{margin-left:0}}.hGxPcf{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1 1 auto;flex:1 1 auto}.tmMkWb{-moz-box-flex:0 1 auto;flex:0 1 auto}.YL9B1{-moz-box-flex:0 0 auto;flex:0 0 auto;margin-top:-0.25rem}.JjRRPc{-moz-box-flex:0 0 auto;flex:0 0 auto;text-align:right}.sMeUxe{margin-right:-1.5rem}.ZjCSDe{margin-top:0.5rem}.jrhqBd.nGmYJe .iCRPId{margin-right:-1rem}.jrhqBd.nGmYJe .WaqnWd,.jrhqBd.nGmYJe .iCRPId{opacity:0.4}.jrhqBd.nGmYJe .cQaDA,.jrhqBd.nGmYJe .tmMkWb,.jrhqBd.nGmYJe .YL9B1,.jrhqBd.nGmYJe .sMeUxe,.jrhqBd.nGmYJe .ZjCSDe,.jrhqBd.nGmYJe .SBOMqf,.jrhqBd.nGmYJe .CEiGpc,.jrhqBd.nGmYJe .YGmIje{opacity:0.67}.CEiGpc,.YGmIje:not(:empty){margin-top:1rem}.x9XmLc .lfGF4,.IGh1ff .lfGF4,.pHPP0b .lfGF4{background-color:#bdc1c6}.x9XmLc .Vlohie,.MejHP .Vlohie,.IGh1ff .Vlohie,.pHPP0b .Vlohie{color:#5f6368}.x9XmLc .tmMkWb,.MejHP .tmMkWb,.IGh1ff .tmMkWb{font-style:italic}.MejHP .tmMkWb{color:#dd2c00}.MejHP .Cm2Nhb{display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;fill:#b31412;margin-right:0.5rem}.n4xnA{padding:0.5rem 0}.DkDwHe{cursor:pointer}.JZicYb{height:3.5rem;padding-right:0.5rem;white-space:nowrap}.qJJSvb{color:#fff;cursor:default;flex-shrink:0;height:2.5rem;line-height:0;margin:0 1rem 0 1.5rem;width:2.5rem}.JZicYb .JRtysb{margin-left:-0.5rem;margin-right:0.5rem}.n8F6Jd{padding:0 1.5rem}.obylVb:not(:empty){margin-bottom:1rem}.rhFKgc{margin-bottom:0.5rem}.s2g3Xd{background-color:transparent;border-top:0.0625rem solid #e0e0e0;overflow:hidden}.JX1kZ[aria-hidden="true"],.ZNE4y:empty{display:none}.ZNE4y{border-top:0.0625rem solid #e0e0e0;box-sizing:border-box;padding:1rem 1.5rem;width:100%}.pablYb{display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;margin:0.5rem 1rem}.GQW44b{overflow:hidden}.tnyRnb{align-self:center;height:2.5rem;margin:0 1rem;width:2.5rem}.tnyRnb:first-child{margin-left:1.5rem}.JEf8lc{flex-shrink:0;margin-right:0.5rem}.qhnNic .UhYXkc{margin-right:1rem;text-align:right}.qhnNic.nGmYJe .qJJSvb,.qhnNic.nGmYJe .JEf8lc{opacity:0.4}.qhnNic.nGmYJe .GQW44b{opacity:0.67}.d4Fe0d{background-color:white;border:0.0625rem solid #dadce0;-moz-border-radius:0.5rem;border-radius:0.5rem;flex-shrink:0;margin-right:1.5rem;padding:1rem;width:10.125rem}.d4Fe0d.s3BYNe{border-color:transparent;padding-top:0;padding-bottom:0}@media (max-width:60rem){.GP1o5c .d4Fe0d{margin-right:0;padding:1rem 1.5rem;width:auto}}@media (max-width:60rem){.zp8Z0e .O0WRkf{background-color:rgba(0,0,0,.12);box-flex:1;flex-grow:1}}.CHJgKd{text-align:right}.uBUej{margin-bottom:-0.5rem;margin-right:-0.5rem}.apFsO{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;display:block}.apFsO.onkcGd,.apFsO.onkcGd:visited{color:rgba(0,0,0,.87)}.oBSRLe{color:rgba(0,0,0,.549);font-weight:500;margin:1rem 0 0 0}.oBSRLe:first-child{margin:0}.sdDCme{color:rgba(0,0,0,.549)}.JwUfNc{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;padding-bottom:.5rem}.oZ63bb{font-weight:500}.hfiB1b{border:0;border-spacing:0}.Gwleff{max-width:10.625rem;padding-right:1rem}.R3OOEd{padding-left:.25rem;padding-right:.25rem}.v9TZ3c{-moz-border-radius:0.5rem;border-radius:0.5rem;margin-top:1.5rem;overflow:hidden}@media (max-width:30em){.v9TZ3c{margin-top:0.5rem}}.qyN25{height:15rem;position:relative;width:100%}.PFLqgc{background-repeat:no-repeat;background-size:cover;height:100%;left:0;position:absolute;top:0;width:100%}@media (max-width:40em){.qyN25{height:11.25rem}}.PFLqgc.KFl4Z:before{background:linear-gradient(rgba(32,33,36,0) 30%,rgba(32,33,36,0.8));content:"";height:100%;left:0;position:absolute;top:0;width:100%}.VVnuU{display:none}.hhj3ub .PFLqgc.PagUde .VVnuU{display:block;height:100%;left:0;opacity:.8;position:absolute;top:0;width:100%}.IzVHde{background-color:#fff;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:space-between}.T4tcpe{bottom:0;color:#fff;left:0;padding:1rem 1.5rem;position:absolute;right:0}@media (max-width:40em){.T4tcpe{padding:1rem 0.5rem}}.T4tcpe.KFl4Z{text-shadow:0 1px 3px rgba(0,0,0,.15),0 1px 2px rgba(0,0,0,.3)}.T4tcpe .tLDEHd{color:#fff}.T4tcpe .tNGpbb,.T4tcpe .qFmcrc{padding-right:2rem}@media (max-width:40em){.T4tcpe .tNGpbb{padding-right:0}}html[dir="rtl"] .PagUde.PFLqgc{transform:scaleX(-1)}.u0Snqb{align-items:center;display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;flex-direction:row}.VkMwfe{margin-right:0.5rem}.uqXhWb.uqXhWb{margin-left:-0.25rem}.VKARh{justify-content:center;bottom:0;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;position:absolute;right:0;width:auto}.lcjGWb{overflow-wrap:break-word}.Y0qupd .v9TZ3c:before{background-image:repeating-linear-gradient(135deg,transparent,transparent 0.5rem,rgba(255,255,255,.3) 0.5rem,rgba(255,255,255,.3) 0.5625rem),repeating-linear-gradient(45deg,rgba(0,0,0,.5),rgba(0,0,0,.5) 0.5rem,rgba(255,255,255,.3) 0.5rem,rgba(255,255,255,.3) 0.5625rem);background-size:0.79549513rem 0.79549513rem;bottom:0;left:0;position:absolute;right:0;top:0}.eZZqMb{position:absolute;right:1rem;top:1rem}.YGy4X{fill:#fff}.GLtrPd{margin-top:0}.NA2Gt{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.NGVAIb{margin-bottom:0.25rem}.RponAc{height:1.5rem;margin-right:0.75rem;width:1.5rem}.MYOkWc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-top:0.5rem}.H0ANOe{width:100%}.UitwCe{margin-top:0.5rem;width:100%}.YiGu3b~.MYOkWc{margin-top:0.25rem}.RHCXAe{margin-left:-0.25rem}.kEAcyb{justify-content:center;margin-top:0.5rem;width:100%}.kEAcyb svg{margin-right:0.25rem}.SDMikc p~p{margin-top:0.5rem}@media not all and (max-width:48.75em){.oT3cQd{display:none}}.QdrXLb[aria-expanded=false] .sTdw3c,.QdrXLb[aria-expanded=true] .JycwX{display:none}.aPHtmf{margin-right:.5rem;display:-moz-inline-box;display:inline-flex;fill:rgb(179,20,18)}.ZK80Pe{padding:0 1.5rem .5rem 0}.ZK80Pe :first-child{-moz-box-flex:1;flex-grow:1}.ZK80Pe .c1OPYd{visibility:hidden}.fcbOGd{flex-shrink:0;margin-right:1rem;width:8rem}.fcbOGd{width:36%}@media (max-width:30rem){.fcbOGd{display:none}}.QdrXLb{margin-bottom:1.5rem}@media (max-width:30rem){.QdrXLb{margin-bottom:1rem}}.QdrXLb:last-child{margin-bottom:0}.G3xBUc{padding:0 1.5rem;position:relative;z-index:0}@media (max-width:30rem){.G3xBUc{padding:0 1rem}}.G3xBUc+.G3xBUc{border-top:.0625rem solid rgb(218,220,224)}@media (max-width:30rem){.c1OPYd{margin-left:1rem}}.OQnryd{display:-moz-box;display:flex;-moz-box-flex:1;flex-grow:1;height:4rem;overflow:hidden}.OQnryd.qwU25c{opacity:1}.OQnryd.qwU25c .UDxXIe{opacity:0.5}.OQnryd.qwU25c .FKELX{opacity:0.27}.UDxXIe{-moz-box-flex:1;flex-grow:1;margin-right:1rem;overflow:hidden}@media (max-width:30rem){.UDxXIe{margin-right:0}}.UDxXIe .SAlC6b{font-weight:500}.vpskfd{-moz-box-flex:1;flex-grow:1;overflow:hidden}@media (max-width:30rem){.vpskfd{display:block}}.vpskfd .IEN71b{color:rgb(213,110,12)}.vpskfd .IEN71b{color:rgb(179,20,18)}.lGVQBf{display:none}@media (max-width:30rem){.lGVQBf{display:block}}.FKELX{margin-right:1rem;color:rgba(0,0,0,.549);line-height:0}.UOYXH{line-height:1;text-align:right}.WMQb5e .oBSRLe{border-top:0.0625rem solid #e0e0e0;padding-top:1rem}.WMQb5e .oBSRLe:first-of-type{border-top:none;padding-top:0}.sxa9Pc{padding-bottom:1rem}.dbEQNc{margin:0 auto;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;width:-moz-calc(100% - 2*1.5rem);width:calc(100% - 2*1.5rem);max-width:62.5rem}.Y0qupd .dbEQNc{max-width:47.5rem}.M7zXZd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-top:1.5rem}.DXLeqd{flex-shrink:0}.Sgw65b{box-flex:1;flex-grow:1}@media not all and (max-width:48.75em){.Sgw65b{overflow:hidden;margin:-1rem;padding:1rem}.rNZeme{display:none}}@media (max-width:48.75em){.DXLeqd .d4Fe0d{margin-right:0;padding:1rem 1.5rem;width:auto}.M7zXZd{flex-direction:column}.dsW6Nd{display:none}}@media (max-width:30em){.dbEQNc{width:auto;flex-direction:column;margin:0 0.5rem}.M7zXZd{margin-top:0.5rem}}.IqBfM{bottom:auto;height:100%;right:auto;width:auto}.vysK6c .dkQQje{display:none}.dkQQje{bottom:1rem;left:1rem;line-height:0;margin:-2px;position:fixed;transition:left .3s cubic-bezier(0,0,0.2,1);z-index:9999}@media (max-width:30em){.dkQQje{bottom:0;left:0}}.QGfKof .dkQQje{left:20.5rem;transition-timing-function:cubic-bezier(0,0,0.2,1)}.OKqsue{z-index:1}.XQOhy>.uyYuVb{left:1.5rem;width:-moz-calc(100% - 1.5rem);width:calc(100% - 1.5rem)}html{overflow:visible}body{overflow:visible;min-height:unset!important}.SSPGKf{min-height:0;height:auto;overflow-y:unset;position:static}.Q001of{bottom:.5rem;color:#333;left:.5rem;position:fixed}.STek2d{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;height:100vh;overflow-x:hidden;overflow-y:auto;position:fixed;z-index:2}.Hlw1k .STek2d{display:none}@media (max-width:65.125rem){.STek2d{display:none}}sentinel{}
/*# sourceURL=/_/mss/boq-apps-edu/_/ss/k=boq-apps-edu.ClassroomUi.TtUpWVPKfDY.L.F4.O/am=BHgWAgAC/d=1/ed=1/rs=AGEDDAsCoucIn376zTYuTYouSXkzYy6Fyg/m=streamview,_b,_tp,_r */</style><script nonce="">onCssLoad();</script><style nonce="">@font-face{font-family:'Roboto';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu72xKOzY.woff2)format('woff2');unicode-range:U+0460-052F,U+1C80-1C88,U+20B4,U+2DE0-2DFF,U+A640-A69F,U+FE2E-FE2F;}@font-face{font-family:'Roboto';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu5mxKOzY.woff2)format('woff2');unicode-range:U+0301,U+0400-045F,U+0490-0491,U+04B0-04B1,U+2116;}@font-face{font-family:'Roboto';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu7mxKOzY.woff2)format('woff2');unicode-range:U+1F00-1FFF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu4WxKOzY.woff2)format('woff2');unicode-range:U+0370-03FF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu7WxKOzY.woff2)format('woff2');unicode-range:U+0102-0103,U+0110-0111,U+0128-0129,U+0168-0169,U+01A0-01A1,U+01AF-01B0,U+1EA0-1EF9,U+20AB;}@font-face{font-family:'Roboto';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu7GxKOzY.woff2)format('woff2');unicode-range:U+0100-024F,U+0259,U+1E00-1EFF,U+2020,U+20A0-20AB,U+20AD-20CF,U+2113,U+2C60-2C7F,U+A720-A7FF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/roboto/v18/KFOmCnqEu92Fr1Mu4mxK.woff2)format('woff2');unicode-range:U+0000-00FF,U+0131,U+0152-0153,U+02BB-02BC,U+02C6,U+02DA,U+02DC,U+2000-206F,U+2074,U+20AC,U+2122,U+2191,U+2193,U+2212,U+2215,U+FEFF,U+FFFD;}@font-face{font-family:'Roboto';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fCRc4EsA.woff2)format('woff2');unicode-range:U+0460-052F,U+1C80-1C88,U+20B4,U+2DE0-2DFF,U+A640-A69F,U+FE2E-FE2F;}@font-face{font-family:'Roboto';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fABc4EsA.woff2)format('woff2');unicode-range:U+0301,U+0400-045F,U+0490-0491,U+04B0-04B1,U+2116;}@font-face{font-family:'Roboto';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fCBc4EsA.woff2)format('woff2');unicode-range:U+1F00-1FFF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fBxc4EsA.woff2)format('woff2');unicode-range:U+0370-03FF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fCxc4EsA.woff2)format('woff2');unicode-range:U+0102-0103,U+0110-0111,U+0128-0129,U+0168-0169,U+01A0-01A1,U+01AF-01B0,U+1EA0-1EF9,U+20AB;}@font-face{font-family:'Roboto';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fChc4EsA.woff2)format('woff2');unicode-range:U+0100-024F,U+0259,U+1E00-1EFF,U+2020,U+20A0-20AB,U+20AD-20CF,U+2113,U+2C60-2C7F,U+A720-A7FF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmEU9fBBc4.woff2)format('woff2');unicode-range:U+0000-00FF,U+0131,U+0152-0153,U+02BB-02BC,U+02C6,U+02DA,U+02DC,U+2000-206F,U+2074,U+20AC,U+2122,U+2191,U+2193,U+2212,U+2215,U+FEFF,U+FFFD;}@font-face{font-family:'Roboto';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfCRc4EsA.woff2)format('woff2');unicode-range:U+0460-052F,U+1C80-1C88,U+20B4,U+2DE0-2DFF,U+A640-A69F,U+FE2E-FE2F;}@font-face{font-family:'Roboto';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfABc4EsA.woff2)format('woff2');unicode-range:U+0301,U+0400-045F,U+0490-0491,U+04B0-04B1,U+2116;}@font-face{font-family:'Roboto';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfCBc4EsA.woff2)format('woff2');unicode-range:U+1F00-1FFF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfBxc4EsA.woff2)format('woff2');unicode-range:U+0370-03FF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfCxc4EsA.woff2)format('woff2');unicode-range:U+0102-0103,U+0110-0111,U+0128-0129,U+0168-0169,U+01A0-01A1,U+01AF-01B0,U+1EA0-1EF9,U+20AB;}@font-face{font-family:'Roboto';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfChc4EsA.woff2)format('woff2');unicode-range:U+0100-024F,U+0259,U+1E00-1EFF,U+2020,U+20A0-20AB,U+20AD-20CF,U+2113,U+2C60-2C7F,U+A720-A7FF;}@font-face{font-family:'Roboto';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/roboto/v18/KFOlCnqEu92Fr1MmWUlfBBc4.woff2)format('woff2');unicode-range:U+0000-00FF,U+0131,U+0152-0153,U+02BB-02BC,U+02C6,U+02DA,U+02DC,U+2000-206F,U+2074,U+20AC,U+2122,U+2191,U+2193,U+2212,U+2215,U+FEFF,U+FFFD;}@font-face{font-family:'Material Icons Extended';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/materialiconsextended/v149/kJEjBvgX7BgnkSrUwT8UnLVc38YydejYY-oE_LvJ.woff2)format('woff2');}.material-icons-extended{font-family:'Material Icons Extended';font-weight:normal;font-style:normal;font-size:24px;line-height:1;letter-spacing:normal;text-transform:none;display:inline-block;white-space:nowrap;word-wrap:normal;direction:ltr;-moz-font-feature-settings:'liga';-moz-osx-font-smoothing:grayscale;}@font-face{font-family:'Google Material Icons';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/googlematerialicons/v130/Gw6kwdfw6UnXLJCcmafZyFRXb3BL9rvi0QZG3Q.woff2)format('woff2');}.google-material-icons{font-family:'Google Material Icons';font-weight:normal;font-style:normal;font-size:24px;line-height:1;letter-spacing:normal;text-transform:none;display:inline-block;white-space:nowrap;word-wrap:normal;direction:ltr;-moz-font-feature-settings:'liga';-moz-osx-font-smoothing:grayscale;}@font-face{font-family:'Product Sans';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/productsans/v9/pxiDypQkot1TnFhsFMOfGShVGdeOcEg.woff2)format('woff2');unicode-range:U+0100-024F,U+0259,U+1E00-1EFF,U+2020,U+20A0-20AB,U+20AD-20CF,U+2113,U+2C60-2C7F,U+A720-A7FF;}@font-face{font-family:'Product Sans';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/productsans/v9/pxiDypQkot1TnFhsFMOfGShVF9eO.woff2)format('woff2');unicode-range:U+0000-00FF,U+0131,U+0152-0153,U+02BB-02BC,U+02C6,U+02DA,U+02DC,U+2000-206F,U+2074,U+20AC,U+2122,U+2191,U+2193,U+2212,U+2215,U+FEFF,U+FFFD;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/googlesans/v14/4UaGrENHsxJlGDuGo1OIlL3Kwp5MKg.woff2)format('woff2');unicode-range:U+0301,U+0400-045F,U+0490-0491,U+04B0-04B1,U+2116;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/googlesans/v14/4UaGrENHsxJlGDuGo1OIlL3Nwp5MKg.woff2)format('woff2');unicode-range:U+0370-03FF;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/googlesans/v14/4UaGrENHsxJlGDuGo1OIlL3Bwp5MKg.woff2)format('woff2');unicode-range:U+0102-0103,U+0110-0111,U+0128-0129,U+0168-0169,U+01A0-01A1,U+01AF-01B0,U+1EA0-1EF9,U+20AB;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/googlesans/v14/4UaGrENHsxJlGDuGo1OIlL3Awp5MKg.woff2)format('woff2');unicode-range:U+0100-024F,U+0259,U+1E00-1EFF,U+2020,U+20A0-20AB,U+20AD-20CF,U+2113,U+2C60-2C7F,U+A720-A7FF;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:400;src:url(//fonts.gstatic.com/s/googlesans/v14/4UaGrENHsxJlGDuGo1OIlL3Owp4.woff2)format('woff2');unicode-range:U+0000-00FF,U+0131,U+0152-0153,U+02BB-02BC,U+02C6,U+02DA,U+02DC,U+2000-206F,U+2074,U+20AC,U+2122,U+2191,U+2193,U+2212,U+2215,U+FEFF,U+FFFD;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLU94Yt3CwZ-Pw.woff2)format('woff2');unicode-range:U+0301,U+0400-045F,U+0490-0491,U+04B0-04B1,U+2116;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLU94YtwCwZ-Pw.woff2)format('woff2');unicode-range:U+0370-03FF;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLU94Yt8CwZ-Pw.woff2)format('woff2');unicode-range:U+0102-0103,U+0110-0111,U+0128-0129,U+0168-0169,U+01A0-01A1,U+01AF-01B0,U+1EA0-1EF9,U+20AB;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLU94Yt9CwZ-Pw.woff2)format('woff2');unicode-range:U+0100-024F,U+0259,U+1E00-1EFF,U+2020,U+20A0-20AB,U+20AD-20CF,U+2113,U+2C60-2C7F,U+A720-A7FF;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:500;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLU94YtzCwY.woff2)format('woff2');unicode-range:U+0000-00FF,U+0131,U+0152-0153,U+02BB-02BC,U+02C6,U+02DA,U+02DC,U+2000-206F,U+2074,U+20AC,U+2122,U+2191,U+2193,U+2212,U+2215,U+FEFF,U+FFFD;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLV154t3CwZ-Pw.woff2)format('woff2');unicode-range:U+0301,U+0400-045F,U+0490-0491,U+04B0-04B1,U+2116;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLV154twCwZ-Pw.woff2)format('woff2');unicode-range:U+0370-03FF;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLV154t8CwZ-Pw.woff2)format('woff2');unicode-range:U+0102-0103,U+0110-0111,U+0128-0129,U+0168-0169,U+01A0-01A1,U+01AF-01B0,U+1EA0-1EF9,U+20AB;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLV154t9CwZ-Pw.woff2)format('woff2');unicode-range:U+0100-024F,U+0259,U+1E00-1EFF,U+2020,U+20A0-20AB,U+20AD-20CF,U+2113,U+2C60-2C7F,U+A720-A7FF;}@font-face{font-family:'Google Sans';font-style:normal;font-weight:700;src:url(//fonts.gstatic.com/s/googlesans/v14/4UabrENHsxJlGDuGo1OIlLV154tzCwY.woff2)format('woff2');unicode-range:U+0000-00FF,U+0131,U+0152-0153,U+02BB-02BC,U+02C6,U+02DA,U+02DC,U+2000-206F,U+2074,U+20AC,U+2122,U+2191,U+2193,U+2212,U+2215,U+FEFF,U+FFFD;}</style><script nonce="">(function(){/*

 Copyright The Closure Library Authors.
 SPDX-License-Identifier: Apache-2.0
*/
'use strict';function aa(){var b=t,c=0;return function(){return c<b.length?{done:!1,value:b[c++]}:{done:!0}}}var w=this||self;/*

 Copyright 2013 Google LLC.
 SPDX-License-Identifier: Apache-2.0
*/
var x={};function ba(b,c){if(null===c)return!1;if("contains"in b&&1==c.nodeType)return b.contains(c);if("compareDocumentPosition"in b)return b==c||!!(b.compareDocumentPosition(c)&16);for(;c&&b!=c;)c=c.parentNode;return c==b};/*

 Copyright 2011 Google LLC.
 SPDX-License-Identifier: Apache-2.0
*/
function ca(b,c){return function(d){d||(d=window.event);return c.call(b,d)}}function y(b){b=b.target||b.srcElement;!b.getAttribute&&b.parentNode&&(b=b.parentNode);return b}var B="undefined"!=typeof navigator&&/Macintosh/.test(navigator.userAgent),da="undefined"!=typeof navigator&&!/Opera/.test(navigator.userAgent)&&/WebKit/.test(navigator.userAgent),ea={A:1,INPUT:1,TEXTAREA:1,SELECT:1,BUTTON:1};function fa(){this._mouseEventsPrevented=!0}
var ha={Enter:13," ":32},C={A:13,BUTTON:0,CHECKBOX:32,COMBOBOX:13,FILE:0,GRIDCELL:13,LINK:13,LISTBOX:13,MENU:0,MENUBAR:0,MENUITEM:0,MENUITEMCHECKBOX:0,MENUITEMRADIO:0,OPTION:0,RADIO:32,RADIOGROUP:32,RESET:0,SUBMIT:0,SWITCH:32,TAB:0,TREE:13,TREEITEM:13},E={CHECKBOX:!0,FILE:!0,OPTION:!0,RADIO:!0},F={COLOR:!0,DATE:!0,DATETIME:!0,"DATETIME-LOCAL":!0,EMAIL:!0,MONTH:!0,NUMBER:!0,PASSWORD:!0,RANGE:!0,SEARCH:!0,TEL:!0,TEXT:!0,TEXTAREA:!0,TIME:!0,URL:!0,WEEK:!0},ia={A:!0,AREA:!0,BUTTON:!0,DIALOG:!0,IMG:!0,
INPUT:!0,LINK:!0,MENU:!0,OPTGROUP:!0,OPTION:!0,PROGRESS:!0,SELECT:!0,TEXTAREA:!0};function ja(b){this.g=b;this.h=[]};var G=w._jsa||{};G._cfc=void 0;G._aeh=void 0;/*

 Copyright 2005 Google LLC.
 SPDX-License-Identifier: Apache-2.0
*/
function L(){this.o=[];this.g=[];this.j=[];this.m={};this.h=null;this.l=[]}function M(b){return String.prototype.trim?b.trim():b.replace(/^\s+/,"").replace(/\s+$/,"")}
function ka(b,c){return function n(a,k){k=void 0===k?!0:k;var e=c;if("click"==e&&(B&&a.metaKey||!B&&a.ctrlKey||2==a.which||null==a.which&&4==a.button||a.shiftKey))e="clickmod";else{var f=a.which||a.keyCode;!f&&a.key&&(f=ha[a.key]);da&&3==f&&(f=13);if(13!=f&&32!=f)f=!1;else{var g=y(a),h;(h="keydown"!=a.type||!!(!("getAttribute"in g)||(g.getAttribute("type")||g.tagName).toUpperCase()in F||"BUTTON"==g.tagName.toUpperCase()||g.type&&"FILE"==g.type.toUpperCase()||g.isContentEditable)||a.ctrlKey||a.shiftKey||
a.altKey||a.metaKey||(g.getAttribute("type")||g.tagName).toUpperCase()in E&&32==f)||((h=g.tagName in ea)||(h=g.getAttributeNode("tabindex"),h=null!=h&&h.specified),h=!(h&&!g.disabled));if(h)f=!1;else{h=(g.getAttribute("role")||g.type||g.tagName).toUpperCase();var v=!(h in C)&&13==f;g="INPUT"!=g.tagName.toUpperCase()||!!g.type;f=(0==C[h]%f||v)&&g}}f&&(e="clickkey")}g=a.srcElement||a.target;f=N(e,a,g,"",null);var l,z;for(h=g;h&&h!=this;h=h.__owner||("#document-fragment"!==(null==(l=h.parentNode)?void 0:
l.nodeName)?h.parentNode:null==(z=h.parentNode)?void 0:z.host)){var m=h;var q=void 0;v=m;var r=e,la=a;var p=v.__jsaction;if(!p){var D;p=null;"getAttribute"in v&&(p=v.getAttribute("jsaction"));if(D=p){p=x[D];if(!p){p={};for(var H=D.split(ma),na=H?H.length:0,I=0;I<na;I++){var A=H[I];if(A){var J=A.indexOf(":"),T=-1!=J;p[T?M(A.substr(0,J)):oa]=T?M(A.substr(J+1)):A}}x[D]=p}v.__jsaction=p}else p=pa,v.__jsaction=p}"maybe_click"==r&&p.click?(q=r,r="click"):"clickkey"==r?r="click":"click"!=r||p.click||(r=
"clickonly");q=G._cfc&&p.click?G._cfc(v,la,p,r,q):{eventType:q?q:r,action:p[r]||"",event:null,ignore:!1};if(q.ignore||q.action)break}q&&(f=N(q.eventType,q.event||a,g,q.action||"",m,f.timeStamp));f&&"touchend"==f.eventType&&(f.event._preventMouseEvents=fa);if(q&&q.action){if(l="clickkey"==e)l=y(a),l=(l.type||l.tagName).toUpperCase(),(l=32==(a.which||a.keyCode)&&"CHECKBOX"!=l)||(l=y(a),z=l.tagName.toUpperCase(),g=(l.getAttribute("role")||"").toUpperCase(),l="BUTTON"===z||"BUTTON"===g?!0:!(l.tagName.toUpperCase()in
ia)||"A"===z||"SELECT"===z||(l.getAttribute("type")||l.tagName).toUpperCase()in E||(l.getAttribute("type")||l.tagName).toUpperCase()in F?!1:!0);l&&(a.preventDefault?a.preventDefault():a.returnValue=!1);if("mouseenter"==e||"mouseleave"==e||"pointerenter"==e||"pointerleave"==e)if(l=a.relatedTarget,!("mouseover"==a.type&&"mouseenter"==e||"mouseout"==a.type&&"mouseleave"==e||"pointerover"==a.type&&"pointerenter"==e||"pointerout"==a.type&&"pointerleave"==e)||l&&(l===m||ba(m,l)))f.action="",f.actionElement=
null;else{e={};for(var u in a)"function"!==typeof a[u]&&"srcElement"!==u&&"target"!==u&&(e[u]=a[u]);e.type="mouseover"==a.type?"mouseenter":"mouseout"==a.type?"mouseleave":"pointerover"==a.type?"pointerenter":"pointerleave";e.target=e.srcElement=m;e.bubbles=!1;f.event=e;f.targetElement=m}}else f.action="",f.actionElement=null;m=f;b.h&&!m.event.a11ysgd&&(u=N(m.eventType,m.event,m.targetElement,m.action,m.actionElement,m.timeStamp),"clickonly"==u.eventType&&(u.eventType="click"),b.h(u,!0));if(m.actionElement){if(b.h){if(!m.actionElement||
"A"!=m.actionElement.tagName||"click"!=m.eventType&&"clickmod"!=m.eventType||(a.preventDefault?a.preventDefault():a.returnValue=!1),(a=b.h(m))&&k){n.call(this,a,!1);return}}else{if((k=w.document)&&!k.createEvent&&k.createEventObject)try{var K=k.createEventObject(a)}catch(ua){K=a}else K=a;m.event=K;b.l.push(m)}G._aeh&&G._aeh(m)}}}function N(b,c,d,a,k,n){return{eventType:b,event:c,targetElement:d,action:a,actionElement:k,timeStamp:n||Date.now()}}
function qa(b,c){return function(d){var a=b,k=c,n=!1;"mouseenter"==a?a="mouseover":"mouseleave"==a?a="mouseout":"pointerenter"==a?a="pointerover":"pointerleave"==a&&(a="pointerout");if(d.addEventListener){if("focus"==a||"blur"==a||"error"==a||"load"==a||"toggle"==a)n=!0;d.addEventListener(a,k,n)}else d.attachEvent&&("focus"==a?a="focusin":"blur"==a&&(a="focusout"),k=ca(d,k),d.attachEvent("on"+a,k));return{eventType:a,i:k,capture:n}}}
function O(b,c,d){if(!b.m.hasOwnProperty(c)){var a=ka(b,c);d=qa(d||c,a);b.m[c]=a;b.o.push(d);for(a=0;a<b.g.length;++a){var k=b.g[a];k.h.push(d.call(null,k.g))}"click"==c&&O(b,"keydown")}}L.prototype.i=function(b){return this.m[b]};
function ra(b,c){var d=new ja(c);a:{for(var a=0;a<b.g.length;a++)if(P(b.g[a].g,c)){c=!0;break a}c=!1}if(c)return b.j.push(d),d;Q(b,d);b.g.push(d);c=b.j.concat(b.g);a=[];for(var k=[],n=0;n<b.g.length;++n){var e=b.g[n];if(R(e,c)){a.push(e);for(var f=0;f<e.h.length;++f){var g=e.g,h=e.h[f];g.removeEventListener?g.removeEventListener(h.eventType,h.i,h.capture):g.detachEvent&&g.detachEvent("on"+h.eventType,h.i)}e.h=[]}else k.push(e)}for(n=0;n<b.j.length;++n)e=b.j[n],R(e,c)?a.push(e):(k.push(e),Q(b,e));
b.g=k;b.j=a;return d}function Q(b,c){var d=c.g;sa&&(d.style.cursor="pointer");for(d=0;d<b.o.length;++d)c.h.push(b.o[d].call(null,c.g))}function R(b,c){for(var d=0;d<c.length;++d)if(c[d].g!=b.g&&P(c[d].g,b.g))return!0;return!1}function P(b,c){for(;b!=c&&c.parentNode;)c=c.parentNode;return b==c}var sa="undefined"!=typeof navigator&&/iPhone|iPad|iPod/.test(navigator.userAgent),ma=/\s*;\s*/,oa="click",pa={};var t="click dblclick focus focusin blur error focusout keydown keyup keypress load mouseover mouseout mouseenter mouseleave submit toggle touchstart touchend touchmove touchcancel auxclick change compositionstart compositionupdate compositionend beforeinput input textinput copy cut paste mousedown mouseup wheel contextmenu dragover dragenter dragleave drop dragstart dragend pointerdown pointermove pointerup pointercancel pointerenter pointerleave pointerover pointerout gotpointercapture lostpointercapture ended loadedmetadata pagehide pageshow visibilitychange beforematch".split(" ");
if(!(t instanceof Array)){var S;var U="undefined"!=typeof Symbol&&Symbol.iterator&&t[Symbol.iterator];if(U)S=U.call(t);else if("number"==typeof t.length)S={next:aa()};else throw Error(String(t)+" is not an iterable or ArrayLike");for(var V,ta=[];!(V=S.next()).done;)ta.push(V.value)};var W=function(b){return{trigger:function(c){var d=b.i(c.type);d||(O(b,c.type),d=b.i(c.type));var a=c.target||c.srcElement;d&&d.call(a.ownerDocument.documentElement,c)},bind:function(c){b.h=c;b.l&&(0<b.l.length&&c(b.l),b.l=null)}}}(function(){var b=window,c=new L,d=ra(c,b.document.documentElement);t.forEach(function(n){return O(c,n)});var a,k;"onwebkitanimationend"in b&&(a="webkitAnimationEnd");O(c,"animationend",a);"onwebkittransitionend"in b&&(k="webkitTransitionEnd");O(c,"transitionend",k);return{s:c,
u:d}}().s),X=["BOQ_wizbind"],Y=window||w;X[0]in Y||"undefined"==typeof Y.execScript||Y.execScript("var "+X[0]);for(var Z;X.length&&(Z=X.shift());)X.length||void 0===W?Y[Z]&&Y[Z]!==Object.prototype[Z]?Y=Y[Z]:Y=Y[Z]={}:Y[Z]=W;}).call(this);
</script><script nocollect="" src="dec2_to_4_files/m=_b,_tp,_r" defer="defer" id="base-js" nonce=""></script><script nonce="">if (window.BOQ_loadedInitialJS) {onJsLoad();} else {document.getElementById('base-js').addEventListener('load', onJsLoad, false);}</script><script nonce="">
    window['_wjdc'] = function (d) {window['_wjdd'] = d};
    </script><style nonce="">.gb_8a:not(.gb_Pd){font:13px/27px Roboto,Arial,sans-serif;z-index:986}@-moz-keyframes gb__a{0%{opacity:0}50%{opacity:1}}@keyframes gb__a{0%{opacity:0}50%{opacity:1}}a.gb_fa{border:none;color:#4285f4;cursor:default;font-weight:bold;outline:none;position:relative;text-align:center;text-decoration:none;text-transform:uppercase;white-space:nowrap;-moz-user-select:none}a.gb_fa:hover:after,a.gb_fa:focus:after{background-color:rgba(0,0,0,.12);content:"";height:100%;left:0;position:absolute;top:0;width:100%}a.gb_fa:hover,a.gb_fa:focus{text-decoration:none}a.gb_fa:active{background-color:rgba(153,153,153,.4);text-decoration:none}a.gb_ga{background-color:#4285f4;color:#fff}a.gb_ga:active{background-color:#0043b2}.gb_ha{-moz-box-shadow:0 1px 1px rgba(0,0,0,.16);box-shadow:0 1px 1px rgba(0,0,0,.16)}.gb_fa,.gb_ga,.gb_ia,.gb_ja{display:inline-block;line-height:28px;padding:0 12px;-moz-border-radius:2px;border-radius:2px}.gb_ia{background:#f8f8f8;border:1px solid #c6c6c6}.gb_ja{background:#f8f8f8}.gb_ia,#gb a.gb_ia.gb_ia,.gb_ja{color:#666;cursor:default;text-decoration:none}#gb a.gb_ja.gb_ja{cursor:default;text-decoration:none}.gb_ja{border:1px solid #4285f4;font-weight:bold;outline:none;background:#4285f4;background:-moz-linear-gradient(top,#4387fd,#4683ea);background:linear-gradient(top,#4387fd,#4683ea);filter:progid:DXImageTransform.Microsoft.gradient(startColorstr=#4387fd,endColorstr=#4683ea,GradientType=0)}#gb a.gb_ja.gb_ja{color:#fff}.gb_ja:hover{-moz-box-shadow:0 1px 0 rgba(0,0,0,.15);box-shadow:0 1px 0 rgba(0,0,0,.15)}.gb_ja:active{-moz-box-shadow:inset 0 2px 0 rgba(0,0,0,.15);box-shadow:inset 0 2px 0 rgba(0,0,0,.15);background:#3c78dc;background:-moz-linear-gradient(top,#3c7ae4,#3f76d3);background:linear-gradient(top,#3c7ae4,#3f76d3);filter:progid:DXImageTransform.Microsoft.gradient(startColorstr=#3c7ae4,endColorstr=#3f76d3,GradientType=0)}#gb .gb_la{background:#fff;border:1px solid #dadce0;color:#1a73e8;display:inline-block;text-decoration:none}#gb .gb_la:hover{background:#f8fbff;border-color:#dadce0;color:#174ea6}#gb .gb_la:focus{background:#f4f8ff;color:#174ea6;outline:1px solid #174ea6}#gb .gb_la:active,#gb .gb_la:focus:active{background:#ecf3fe;color:#174ea6}#gb .gb_la.gb_g{background:transparent;border:1px solid #5f6368;color:#8ab4f8;text-decoration:none}#gb .gb_la.gb_g:hover{background:rgba(255,255,255,.04);color:#e8eaed}#gb .gb_la.gb_g:focus{background:rgba(232,234,237,.12);color:#e8eaed;outline:1px solid #e8eaed}#gb .gb_la.gb_g:active,#gb .gb_la.gb_g:focus:active{background:rgba(232,234,237,.1);color:#e8eaed}.gb_j{display:none!important}.gb_Ra{visibility:hidden}.gb_od{display:inline-block;vertical-align:middle}.gb_Ef .gb_i{bottom:-3px;right:-5px}.gb_Ff{position:relative}.gb_e{display:inline-block;outline:none;vertical-align:middle;-moz-border-radius:2px;border-radius:2px;-moz-box-sizing:border-box;box-sizing:border-box;height:40px;width:40px;color:#000;cursor:pointer;text-decoration:none}#gb#gb a.gb_e{color:#000;cursor:pointer;text-decoration:none}.gb_ab{border-color:transparent;border-bottom-color:#fff;border-style:dashed dashed solid;border-width:0 8.5px 8.5px;display:none;position:absolute;left:11.5px;top:43px;z-index:1;height:0;width:0;-moz-animation:gb__a .2s;animation:gb__a .2s}.gb_bb{border-color:transparent;border-style:dashed dashed solid;border-width:0 8.5px 8.5px;display:none;position:absolute;left:11.5px;z-index:1;height:0;width:0;-moz-animation:gb__a .2s;animation:gb__a .2s;border-bottom-color:#ccc;border-bottom-color:rgba(0,0,0,.2);top:42px}x:-o-prefocus,div.gb_bb{border-bottom-color:#ccc}.gb_P{background:#fff;border:1px solid #ccc;border-color:rgba(0,0,0,.2);color:#000;-moz-box-shadow:0 2px 10px rgba(0,0,0,.2);box-shadow:0 2px 10px rgba(0,0,0,.2);display:none;outline:none;overflow:hidden;position:absolute;right:8px;top:62px;-moz-animation:gb__a .2s;animation:gb__a .2s;-moz-border-radius:2px;border-radius:2px;-moz-user-select:text}.gb_od.gb_Ba .gb_ab,.gb_od.gb_Ba .gb_bb,.gb_od.gb_Ba .gb_P,.gb_Ba.gb_P{display:block}.gb_od.gb_Ba.gb_Hf .gb_ab,.gb_od.gb_Ba.gb_Hf .gb_bb{display:none}.gb_If{position:absolute;right:8px;top:62px;z-index:-1}.gb_Xa .gb_ab,.gb_Xa .gb_bb,.gb_Xa .gb_P{margin-top:-10px}.gb_od:first-child,#gbsfw:first-child+.gb_od{padding-left:4px}.gb_Fa.gb_We .gb_od:first-child{padding-left:0}.gb_Xe{position:relative}.gb_0c .gb_Xe,.gb_6d .gb_Xe{float:right}.gb_e{padding:8px;cursor:pointer}.gb_Fa .gb_gd:not(.gb_fa):focus img{background-color:rgba(0,0,0,.20);outline:none;-moz-border-radius:50%;border-radius:50%}.gb_Ze button svg,.gb_e{-moz-border-radius:50%;border-radius:50%}.gb_Ze button:focus:not(:focus-visible) svg,.gb_Ze button:hover svg,.gb_Ze button:active svg,.gb_e:focus:not(:focus-visible),.gb_e:hover,.gb_e:active,.gb_e[aria-expanded=true]{outline:none}.gb_Jc .gb_Ze.gb_0e button:focus-visible svg,.gb_Ze button:focus-visible svg,.gb_e:focus-visible{outline:1px solid #202124}.gb_Jc .gb_Ze button:focus-visible svg,.gb_Jc .gb_e:focus-visible{outline:1px solid #f1f3f4}@media (forced-colors:active){.gb_Jc .gb_Ze.gb_0e button:focus-visible svg,.gb_Ze button:focus-visible svg,.gb_Jc .gb_Ze button:focus-visible svg{outline:1px solid currentcolor}}.gb_Jc .gb_Ze.gb_0e button:focus svg,.gb_Jc .gb_Ze.gb_0e button:focus:hover svg,.gb_Ze button:focus svg,.gb_Ze button:focus:hover svg,.gb_e:focus,.gb_e:focus:hover{background-color:rgba(60,64,67,.1)}.gb_Jc .gb_Ze.gb_0e button:active svg,.gb_Ze button:active svg,.gb_e:active{background-color:rgba(60,64,67,.12)}.gb_Jc .gb_Ze.gb_0e button:hover svg,.gb_Ze button:hover svg,.gb_e:hover{background-color:rgba(60,64,67,.08)}.gb_za .gb_e.gb_1a:hover{background-color:transparent}.gb_e[aria-expanded=true],.gb_e:hover[aria-expanded=true]{background-color:rgba(95,99,104,.24)}.gb_e[aria-expanded=true] .gb_1e,.gb_e[aria-expanded=true] .gb_2e{fill:#5f6368;opacity:1}.gb_Jc .gb_Ze button:hover svg,.gb_Jc .gb_e:hover{background-color:rgba(232,234,237,.08)}.gb_Jc .gb_Ze button:focus svg,.gb_Jc .gb_Ze button:focus:hover svg,.gb_Jc .gb_e:focus,.gb_Jc .gb_e:focus:hover{background-color:rgba(232,234,237,.10)}.gb_Jc .gb_Ze button:active svg,.gb_Jc .gb_e:active{background-color:rgba(232,234,237,.12)}.gb_Jc .gb_e[aria-expanded=true],.gb_Jc .gb_e:hover[aria-expanded=true]{background-color:rgba(255,255,255,.12)}.gb_Jc .gb_e[aria-expanded=true] .gb_1e,.gb_Jc .gb_e[aria-expanded=true] .gb_2e{fill:#fff;opacity:1}.gb_od{padding:4px}.gb_Fa.gb_We .gb_od{padding:4px 2px}.gb_Fa.gb_We .gb_b.gb_od{padding-left:6px}.gb_P{z-index:991;line-height:normal}.gb_P.gb_3e{left:8px;right:auto}@media (max-width:350px){.gb_P.gb_3e{left:0}}.gb_4e .gb_P{top:56px}.gb_N .gb_e,.gb_O .gb_N .gb_e{background-position:-64px -29px}.gb_t .gb_N .gb_e{background-position:-29px -29px;opacity:1}.gb_N .gb_e,.gb_N .gb_e:hover,.gb_N .gb_e:focus{opacity:1}.gb_Qd{display:none}.gb_i{display:none}.gb_8c{font-family:Google Sans,Roboto,Helvetica,Arial,sans-serif;font-size:20px;font-weight:400;letter-spacing:0.25px;line-height:48px;margin-bottom:2px;opacity:1;overflow:hidden;padding-left:16px;position:relative;text-overflow:ellipsis;vertical-align:middle;top:2px;white-space:nowrap;flex:1 1 auto}.gb_8c.gb_9c{color:#3c4043}.gb_Fa.gb_Ha .gb_8c{margin-bottom:0}.gb_ad.gb_bd .gb_8c{padding-left:4px}.gb_Fa.gb_Ha .gb_cd{position:relative;top:-2px}.gb_Fa{color:black;min-width:320px;position:relative;-moz-transition:box-shadow 250ms;transition:box-shadow 250ms}.gb_Fa.gb_Rc{min-width:240px}.gb_Fa.gb_Rd .gb_Sd{display:none}.gb_Fa.gb_Rd .gb_Td{height:56px}header.gb_Fa{display:block}.gb_Fa svg{fill:currentColor}.gb_Ud{position:fixed;top:0;width:100%}.gb_Vd{-moz-box-shadow:0px 4px 5px 0px rgba(0,0,0,.14),0px 1px 10px 0px rgba(0,0,0,.12),0px 2px 4px -1px rgba(0,0,0,.2);box-shadow:0px 4px 5px 0px rgba(0,0,0,.14),0px 1px 10px 0px rgba(0,0,0,.12),0px 2px 4px -1px rgba(0,0,0,.2)}.gb_Wd{height:64px}.gb_Td{box-sizing:border-box;position:relative;width:100%;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;justify-content:space-between;min-width:-webkit-min-content;min-width:-moz-min-content;min-width:-ms-min-content;min-width:min-content}.gb_Fa:not(.gb_Ha) .gb_Td{padding:8px}.gb_Fa.gb_Xd .gb_Td{flex:1 0 auto}.gb_Fa .gb_Td.gb_Zd.gb_0d{min-width:0}.gb_Fa.gb_Ha .gb_Td{padding:4px;padding-left:8px;min-width:0}.gb_Sd{height:48px;vertical-align:middle;white-space:nowrap;-moz-box-align:center;align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-user-select:-moz-none}.gb_2d>.gb_Sd{display:table-cell;width:100%}.gb_ad{padding-right:30px;-moz-box-sizing:border-box;box-sizing:border-box;flex:1 0 auto}.gb_Fa.gb_Ha .gb_ad{padding-right:14px}.gb_3d{flex:1 1 100%}.gb_3d>:only-child{display:inline-block}.gb_4d.gb_1c{padding-left:4px}.gb_4d.gb_5d,.gb_Fa.gb_Xd .gb_4d,.gb_Fa.gb_Ha:not(.gb_6d) .gb_4d{padding-left:0}.gb_Fa.gb_Ha .gb_4d.gb_5d{padding-right:0}.gb_Fa.gb_Ha .gb_4d.gb_5d .gb_za{margin-left:10px}.gb_1c{display:inline}.gb_Fa.gb_Uc .gb_4d.gb_7d,.gb_Fa.gb_6d .gb_4d.gb_7d{padding-left:2px}.gb_8c{display:inline-block}.gb_4d{box-sizing:border-box;height:48px;line-height:normal;padding:0 4px;padding-left:30px;flex:0 0 auto;justify-content:flex-end}.gb_6d{height:48px}.gb_Fa.gb_6d{min-width:initial;min-width:auto}.gb_6d .gb_4d{float:right;padding-left:32px}.gb_6d .gb_4d.gb_8d{padding-left:0}.gb_9d{font-size:14px;max-width:200px;overflow:hidden;padding:0 12px;text-overflow:ellipsis;white-space:nowrap;-moz-user-select:text}.gb_ae{transition:background-color .4s}.gb_be{color:black}.gb_Jc{color:white}.gb_Fa a,.gb_Oc a{color:inherit}.gb_D{color:rgba(0,0,0,.87)}.gb_Fa svg,.gb_Oc svg,.gb_ad .gb_ce,.gb_0c .gb_ce{color:#5f6368;opacity:1}.gb_Jc svg,.gb_Oc.gb_Sc svg,.gb_Jc .gb_ad .gb_ce,.gb_Jc .gb_ad .gb_Ic,.gb_Jc .gb_ad .gb_cd,.gb_Oc.gb_Sc .gb_ce{color:rgba(255,255,255,0.87)}.gb_Jc .gb_ad .gb_Hc:not(.gb_de){opacity:0.87}.gb_9c{color:inherit;opacity:1;text-rendering:optimizeLegibility;-moz-osx-font-smoothing:grayscale}.gb_Jc .gb_9c,.gb_be .gb_9c{opacity:1}.gb_ee{position:relative}.gb_fe{font-family:arial,sans-serif;line-height:normal;padding-right:15px}a.gb_q,span.gb_q{color:rgba(0,0,0,.87);text-decoration:none}.gb_Jc a.gb_q,.gb_Jc span.gb_q{color:white}a.gb_q:focus{outline-offset:2px}a.gb_q:hover{text-decoration:underline}.gb_r{display:inline-block;padding-left:15px}.gb_r .gb_q{display:inline-block;line-height:24px;vertical-align:middle}.gb_ge{font-family:Google Sans,Roboto,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;letter-spacing:0.25px;line-height:16px;margin-left:10px;margin-right:8px;min-width:96px;padding:9px 23px;text-align:center;vertical-align:middle;-moz-border-radius:4px;border-radius:4px;-moz-box-sizing:border-box;box-sizing:border-box}.gb_Fa.gb_6d .gb_ge{margin-left:8px}#gb a.gb_ja.gb_ja.gb_ge{cursor:pointer}.gb_ja.gb_ge:hover{background:#1b66c9;-moz-box-shadow:0 1px 3px 1px rgba(66,64,67,.15),0 1px 2px 0 rgba(60,64,67,.3);box-shadow:0 1px 3px 1px rgba(66,64,67,.15),0 1px 2px 0 rgba(60,64,67,.3)}.gb_ja.gb_ge:focus,.gb_ja.gb_ge:hover:focus{background:#1c5fba;-moz-box-shadow:0 1px 3px 1px rgba(66,64,67,.15),0 1px 2px 0 rgba(60,64,67,.3);box-shadow:0 1px 3px 1px rgba(66,64,67,.15),0 1px 2px 0 rgba(60,64,67,.3)}.gb_ja.gb_ge:active{background:#1b63c1;-moz-box-shadow:0 1px 3px 1px rgba(66,64,67,.15),0 1px 2px 0 rgba(60,64,67,.3);box-shadow:0 1px 3px 1px rgba(66,64,67,.15),0 1px 2px 0 rgba(60,64,67,.3)}.gb_ge{background:#1a73e8;border:1px solid transparent}.gb_Fa.gb_Ha .gb_ge{padding:9px 15px;min-width:80px}.gb_he{text-align:left}#gb .gb_Jc a.gb_ge:not(.gb_g),#gb.gb_Jc a.gb_ge{background:#fff;border-color:#dadce0;-moz-box-shadow:none;box-shadow:none;color:#1a73e8}#gb a.gb_ja.gb_g.gb_ge{background:#8ab4f8;border:1px solid transparent;-moz-box-shadow:none;box-shadow:none;color:#202124}#gb .gb_Jc a.gb_ge:hover:not(.gb_g),#gb.gb_Jc a.gb_ge:hover{background:#f8fbff;border-color:#cce0fc}#gb a.gb_ja.gb_g.gb_ge:hover{background:#93baf9;border-color:transparent;-moz-box-shadow:0 1px 3px 1px rgba(0,0,0,.15),0 1px 2px rgba(0,0,0,.3);box-shadow:0 1px 3px 1px rgba(0,0,0,.15),0 1px 2px rgba(0,0,0,.3)}#gb .gb_Jc a.gb_ge:focus:not(.gb_g),#gb .gb_Jc a.gb_ge:focus:hover:not(.gb_g),#gb.gb_Jc a.gb_ge:focus:not(.gb_g),#gb.gb_Jc a.gb_ge:focus:hover:not(.gb_g){background:#f4f8ff;outline:1px solid #c9ddfc}#gb a.gb_ja.gb_g.gb_ge:focus,#gb a.gb_ja.gb_g.gb_ge:focus:hover{background:#a6c6fa;border-color:transparent;-moz-box-shadow:none;box-shadow:none}#gb .gb_Jc a.gb_ge:active:not(.gb_g),#gb.gb_Jc a.gb_ge:active{background:#ecf3fe}#gb a.gb_ja.gb_g.gb_ge:active{background:#a1c3f9;-moz-box-shadow:0 1px 2px rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);box-shadow:0 1px 2px rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15)}.gb_za{background-color:rgba(255,255,255,.88);border:1px solid #dadce0;box-sizing:border-box;cursor:pointer;display:inline-block;max-height:48px;overflow:hidden;outline:none;padding:0;vertical-align:middle;width:134px;-moz-border-radius:8px;border-radius:8px}.gb_za.gb_g{background-color:transparent;border:1px solid #5f6368}.gb_Aa{display:inherit}.gb_za.gb_g .gb_Aa{background:#fff;-moz-border-radius:4px;border-radius:4px;display:inline-block;left:8px;margin-right:5px;position:relative;padding:3px;top:-1px}.gb_za:hover{border:1px solid #d2e3fc;background-color:rgba(248,250,255,.88)}.gb_za.gb_g:hover{background-color:rgba(241,243,244,.04);border:1px solid #5f6368}.gb_za:focus-visible,.gb_za:focus{background-color:rgba(255,255,255);outline:1px solid #202124;-moz-box-shadow:0px 1px 2px 0px rgba(60,64,67,.3),0px 1px 3px 1px rgba(60,64,67,.15);box-shadow:0px 1px 2px 0px rgba(60,64,67,.3),0px 1px 3px 1px rgba(60,64,67,.15)}.gb_za.gb_g:focus-visible,.gb_za.gb_g:focus{background-color:rgba(241,243,244,.12);outline:1px solid #f1f3f4;-moz-box-shadow:0 1px 3px 1px rgba(0,0,0,.15),0 1px 2px 0 rgba(0,0,0,.3);box-shadow:0 1px 3px 1px rgba(0,0,0,.15),0 1px 2px 0 rgba(0,0,0,.3)}.gb_za.gb_g:active,.gb_za.gb_Ba.gb_g:focus{background-color:rgba(241,243,244,.1);border:1px solid #5f6368}.gb_Ca{display:inline-block;padding-bottom:2px;padding-left:7px;padding-top:2px;text-align:center;vertical-align:middle;line-height:32px;width:78px}.gb_za.gb_g .gb_Ca{line-height:26px;margin-left:0;padding-bottom:0;padding-left:0;padding-top:0;width:72px}.gb_Ca.gb_Da{background-color:#f1f3f4;-moz-border-radius:4px;border-radius:4px;margin-left:8px;padding-left:0}.gb_Ca.gb_Da .gb_Ea{vertical-align:middle}.gb_Fa:not(.gb_Ha) .gb_za{margin-left:10px;margin-right:4px}.gb_Ia{max-height:32px;width:78px}.gb_za.gb_g .gb_Ia{max-height:26px;width:72px}.gb_h{background-size:32px 32px;border:0;-moz-border-radius:50%;border-radius:50%;display:block;margin:0px;position:relative;height:32px;width:32px;z-index:0}.gb_Sa{background-color:#e8f0fe;border:1px solid rgba(32,33,36,.08);position:relative}.gb_Sa.gb_h{height:30px;width:30px}.gb_Sa.gb_h:hover,.gb_Sa.gb_h:active{-moz-box-shadow:none;box-shadow:none}.gb_Ta{background:#fff;border:none;-moz-border-radius:50%;border-radius:50%;bottom:2px;-moz-box-shadow:0px 1px 2px 0px rgba(60,64,67,.30),0px 1px 3px 1px rgba(60,64,67,.15);box-shadow:0px 1px 2px 0px rgba(60,64,67,.30),0px 1px 3px 1px rgba(60,64,67,.15);height:14px;margin:2px;position:absolute;right:0;width:14px}.gb_Ua{color:#1f71e7;font:400 22px/32px Google Sans,Roboto,Helvetica,Arial,sans-serif;text-align:center;text-transform:uppercase}@media (min-resolution:1.25dppx),(-o-min-device-pixel-ratio:5/4),(-webkit-min-device-pixel-ratio:1.25),(min-device-pixel-ratio:1.25){.gb_h::before,.gb_Va::before{display:inline-block;-moz-transform:scale(.5);transform:scale(.5);-moz-transform-origin:left 0;transform-origin:left 0}.gb_v .gb_Va::before{-moz-transform:scale(0.416666667);transform:scale(0.416666667)}}.gb_h:hover,.gb_h:focus{-moz-box-shadow:0 1px 0 rgba(0,0,0,.15);box-shadow:0 1px 0 rgba(0,0,0,.15)}.gb_h:active{-moz-box-shadow:inset 0 2px 0 rgba(0,0,0,.15);box-shadow:inset 0 2px 0 rgba(0,0,0,.15)}.gb_h:active::after{background:rgba(0,0,0,.1);-moz-border-radius:50%;border-radius:50%;content:"";display:block;height:100%}.gb_Wa{cursor:pointer;line-height:40px;min-width:30px;opacity:.75;overflow:hidden;vertical-align:middle;text-overflow:ellipsis}.gb_e.gb_Wa{width:auto}.gb_Wa:hover,.gb_Wa:focus{opacity:.85}.gb_Xa .gb_Wa,.gb_Xa .gb_Za{line-height:26px}#gb#gb.gb_Xa a.gb_Wa,.gb_Xa .gb_Za{font-size:11px;height:auto}.gb_0a{border-top:4px solid #000;border-left:4px dashed transparent;border-right:4px dashed transparent;display:inline-block;margin-left:6px;opacity:.75;vertical-align:middle}.gb_1a:hover .gb_0a{opacity:.85}.gb_za>.gb_b{padding:3px 3px 3px 4px}.gb_2a.gb_Ra{color:#fff}.gb_t .gb_Wa,.gb_t .gb_0a{opacity:1}#gb#gb.gb_t.gb_t a.gb_Wa,#gb#gb .gb_t.gb_t a.gb_Wa{color:#fff}.gb_t.gb_t .gb_0a{border-top-color:#fff;opacity:1}.gb_O .gb_h:hover,.gb_t .gb_h:hover,.gb_O .gb_h:focus,.gb_t .gb_h:focus{-moz-box-shadow:0 1px 0 rgba(0,0,0,.15),0 1px 2px rgba(0,0,0,.2);box-shadow:0 1px 0 rgba(0,0,0,.15),0 1px 2px rgba(0,0,0,.2)}.gb_3a .gb_b,.gb_4a .gb_b{position:absolute;right:1px}.gb_b.gb_s,.gb_5a.gb_s,.gb_1a.gb_s{flex:0 1 auto;flex:0 1 main-size}.gb_6a.gb_7a .gb_Wa{width:30px!important}.gb_d{height:40px;position:absolute;right:-5px;top:-5px;width:40px}.gb_8a .gb_d,.gb_9a .gb_d{right:0;top:0}.gb_b .gb_e{padding:4px}.gb_k{display:none}sentinel{}</style><script nonce="">;this.gbar_={CONFIG:[[[0,"www.gstatic.com","og.qtm.en_US.ODCNLawGeLk.2019.O","com.br","pt-BR","265",0,[4,2,"","","","517837492","0"],null,"ShkiZMnGFf-GwbkPztue2AE",null,0,"og.qtm._w-zyUPsPZw.L.F4.O","AA2YrTvkbJWV1adPbuzYq0DsgPYnetf7Bg","AA2YrTvmtKM57xcbKdJeX3djH0NMhQr_Nw","",2,1,200,"BRA",null,null,"269","265",1],null,[1,0.1000000014901161,2,1],[1,0.001000000047497451,1],[1,0,1,null,"0","r243360@dac.unicamp.br","","AEq3ON3Glse3dF_KXFnOaewsCdQHwMtF0ajoX5d1tDmA1yMLx8LVVZZAIeUx19I0tq6-EKeyOCW9sYp2PrTjO9FWDWEaj3YCiQ"],[0,0,"",1,0,0,0,0,0,0,null,0,0,null,0,0,null,null,0,0,0,"","","","","","",null,0,0,0,0,0,null,null,null,"rgba(32,33,36,1)","rgba(255,255,255,1)",0,0,1,null,null,1,0,0],["%1$s (padrão)","Conta de marca",1,"%1$s (delegada)",1,null,83,"/c/NDQ4MTYxOTM2MzI4?authuser=$authuser",null,null,null,1,"https://accounts.google.com/ListAccounts?authuser=0\u0026pid=265\u0026gpsia=1\u0026source=ogb\u0026atic=1\u0026mo=1\u0026mn=1\u0026hl=pt-BR\u0026ts=102",0,"dashboard",null,null,null,null,"Perfil","",1,null,"Desconectada","https://accounts.google.com/AccountChooser?source=ogb\u0026continue=$continue\u0026Email=$email\u0026ec=GAhAiQI","https://accounts.google.com/RemoveLocalAccount?source=ogb","Remover","Fazer login",0,1,1,0,1,1,0,null,null,null,"Sessão expirada",null,null,null,"Visitante",null,"Padrão","Delegada","Sair de todas as contas",1,null,null,0,null,null,"myaccount.google.com","https",0,1,0],null,["1","gci_91f30755d6a6b787dcc2a4062e6e9824.js","googleapis.client:gapi.iframes","0","pt-BR"],null,null,null,null,["m;/_/scs/abc-static/_/js/k=gapi.gapi.en.fpEXMBCWMKc.O/d=1/rs=AHpOoo9SQGHwxhl93I-W5KEIEdf87vGuqQ/m=__features__","https://apis.google.com","","","1","",null,1,"es_plusone_gc_20230306.0_p1","pt-BR",null,0],[0.009999999776482582,"com.br","265",[null,"","0",null,1,5184000,null,null,"",null,null,null,null,null,0,null,0,0,1,0,0,0,null,null,0,0,null,0,0,0,0,0],null,null,null,0,null,null,["5061451","google\\.(com|ru|ca|by|kz|com\\.mx|com\\.tr)$",1]],[1,1,null,40400,265,"BRA","pt-BR","517837492.0",8,0.009999999776482582,1,0,null,null,null,null,"3701102,3701113,3701124",null,null,null,"ShkiZMnGFf-GwbkPztue2AE",0,0,0,null,2,5,"ug",119,0,0,1,0,1],[[null,null,null,"https://www.gstatic.com/og/_/js/k=og.qtm.en_US.ODCNLawGeLk.2019.O/rt=j/m=qabr,qgl,q_dnp,qcwid,qbd,qapid,qrcd/exm=qaaw,qadd,qaid,qein,qhaw,qhba,qhbr,qhch,qhga,qhid,qhin,qhpr/d=1/ed=1/rs=AA2YrTvkbJWV1adPbuzYq0DsgPYnetf7Bg"],[null,null,null,"https://www.gstatic.com/og/_/ss/k=og.qtm._w-zyUPsPZw.L.F4.O/m=qcwid/excm=qaaw,qadd,qaid,qein,qhaw,qhba,qhbr,qhch,qhga,qhid,qhin,qhpr/d=1/ed=1/ct=zgms/rs=AA2YrTvmtKM57xcbKdJeX3djH0NMhQr_Nw"]],null,null,null,[[[null,null,[null,null,null,"https://ogs.google.com/u/0/widget/app?awv2=1"],0,448,328,57,4,1,0,0,63,64,8000,"https://www.google.com.br/intl/pt-BR/about/products",67,1,69,null,1,70,"Ocorreu um problema no carregamento do conjunto de aplicativos. Tente novamente em alguns minutos ou acesse a página %1$sProdutos do Google%2$s.",3,0,0,74,4000,null,null,null,null,null,null,null,"/widget/app",null,null,null,null,null,null,null,0],[null,null,[null,null,null,"https://ogs.google.com/u/0/widget/account?amf=1\u0026sea=1"],0,414,400,57,4,1,0,0,65,66,8000,"https://accounts.google.com/SignOutOptions?hl=pt-BR\u0026continue=https://classroom.google.com/c/NDQ4MTYxOTM2MzI4",68,2,null,null,1,113,"Algo deu errado. Atualize para tentar novamente ou %1$sescolha outra conta%2$s.",3,null,null,75,0,null,null,null,null,null,null,null,"/widget/account",["https","myaccount.google.com",0,32,83,0],0,0,1,["Alerta crítico de segurança","Alerta importante da conta"],0,1,0]],null,null,"269","265",1,0,null,"pt-BR",0,["/c/NDQ4MTYxOTM2MzI4?authuser=$authuser","https://accounts.google.com/AddSession?service=classroom\u0026continue=https://classroom.google.com/c/NDQ4MTYxOTM2MzI4\u0026ec=GAlAiQI","https://accounts.google.com/Logout?ec=GAdAiQI","https://accounts.google.com/ListAccounts?authuser=0\u0026pid=265\u0026gpsia=1\u0026source=ogb\u0026atic=1\u0026mo=1\u0026mn=1\u0026hl=pt-BR\u0026ts=102",0,0,"",0,0,null,0,0],0,0,0,null,0],null,[["mousedown","touchstart","touchmove","wheel","keydown"],300000],[[null,null,null,"https://accounts.google.com/RotateCookiesPage"],3,4000,1]]],};this.gbar_=this.gbar_||{};(function(_){var window=this;
try{
/*

 Copyright The Closure Library Authors.
 SPDX-License-Identifier: Apache-2.0
*/
var ta,Ja,Ka,La,Na,Ta,Va,Ua,Xa,Ya,Za,cb,$a,fb,gb;_.ba=function(a,b){if(Error.captureStackTrace)Error.captureStackTrace(this,_.ba);else{const c=Error().stack;c&&(this.stack=c)}a&&(this.message=String(a));void 0!==b&&(this.cause=b)};_.ca=function(){var a=_.m.navigator;return a&&(a=a.userAgent)?a:""};_.fa=function(a){return da?_.ea?_.ea.brands.some(({brand:b})=>b&&-1!=b.indexOf(a)):!1:!1};_.n=function(a){return-1!=_.ca().indexOf(a)};_.ha=function(){return da?!!_.ea&&0<_.ea.brands.length:!1};
_.ia=function(){return _.ha()?!1:_.n("Opera")};_.ja=function(){return _.ha()?!1:_.n("Trident")||_.n("MSIE")};_.ka=function(){return _.ha()?!1:_.n("Edge")};_.la=function(){return _.ha()?_.fa("Microsoft Edge"):_.n("Edg/")};_.ma=function(){return _.n("Firefox")||_.n("FxiOS")};_.oa=function(){return _.n("Safari")&&!(_.na()||(_.ha()?0:_.n("Coast"))||_.ia()||_.ka()||_.la()||(_.ha()?_.fa("Opera"):_.n("OPR"))||_.ma()||_.n("Silk")||_.n("Android"))};
_.na=function(){return _.ha()?_.fa("Chromium"):(_.n("Chrome")||_.n("CriOS"))&&!_.ka()||_.n("Silk")};_.pa=function(){return _.n("Android")&&!(_.na()||_.ma()||_.ia()||_.n("Silk"))};_.ra=function(){return da?!!_.ea&&!!_.ea.platform:!1};_.sa=function(){return _.ra()?"Android"===_.ea.platform:_.n("Android")};ta=function(){return _.n("iPhone")&&!_.n("iPod")&&!_.n("iPad")};_.ua=function(){return ta()||_.n("iPad")||_.n("iPod")};_.va=function(){return _.ra()?"macOS"===_.ea.platform:_.n("Macintosh")};
_.wa=function(){return _.ra()?"Windows"===_.ea.platform:_.n("Windows")};_.xa=function(a){const b=a.length;if(0<b){const c=Array(b);for(let d=0;d<b;d++)c[d]=a[d];return c}return[]};_.ya=function(){return-1!=_.ca().toLowerCase().indexOf("webkit")&&!_.n("Edge")};_.Ba=function(a){if(!_.za)return _.Aa(a);let b="";for(;10240<a.length;)b+=String.fromCharCode.apply(null,a.subarray(0,10240)),a=a.subarray(10240);b+=String.fromCharCode.apply(null,a);return btoa(b)};
_.Da=function(a){return Ca&&null!=a&&a instanceof Uint8Array};_.Fa=function(a,b){if(_.Ea)return a[_.Ea]|=b;if(void 0!==a.Bb)return a.Bb|=b;Object.defineProperties(a,{Bb:{value:b,configurable:!0,writable:!0,enumerable:!1}});return b};_.r=function(a){let b;_.Ea?b=a[_.Ea]:b=a.Bb;return null==b?0:b};_.Ga=function(a,b){_.Ea?a[_.Ea]=b:void 0!==a.Bb?a.Bb=b:Object.defineProperties(a,{Bb:{value:b,configurable:!0,writable:!0,enumerable:!1}});return a};_.Ha=function(a){_.Fa(a,1);return a};
_.Ia=function(a){_.Fa(a,16);return a};Ja=function(a,b){_.Ga(b,(a|0)&-51)};Ka=function(a,b){_.Ga(b,(a|18)&-41)};La=function(a){return null!==a&&"object"===typeof a&&!Array.isArray(a)&&a.constructor===Object};_.Ma=function(a){if(_.r(a.na)&2)throw Error();};Na=function(a){var b=a.length;(b=b?a[b-1]:void 0)&&La(b)?b.g=1:a.push({g:1})};_.Oa=function(a,b){const c=_.r(a);let d=c;0===d&&(d|=b&16);d|=b&2;d!==c&&_.Ga(a,d)};_.Pa=function(a,b){return null==a?b:a};
_.Ra=function(a,b){Qa=b;a=new a(b);Qa=void 0;return a};Ta=function(a){switch(typeof a){case "number":return isFinite(a)?a:String(a);case "object":if(a)if(Array.isArray(a)){if(0!==(_.r(a)&128))return a=Array.prototype.slice.call(a),Na(a),a}else{if(_.Da(a))return _.Ba(a);if("function"==typeof _.Sa&&a instanceof _.Sa)return a.j()}}return a};
Va=function(a,b,c,d,e){if(null!=a){if(Array.isArray(a))a=e&&0==a.length&&_.r(a)&1?void 0:Ua(a,b,c,void 0!==d,e);else if(La(a)){const f={};for(let g in a)f[g]=Va(a[g],b,c,d,e);a=f}else a=b(a,d);return a}};Ua=function(a,b,c,d,e){const f=_.r(a);d=d?!!(f&16):void 0;a=Array.prototype.slice.call(a);for(let g=0;g<a.length;g++)a[g]=Va(a[g],b,c,d,e);c(f,a);return a};Xa=function(a){return a.ie===Wa?a.toJSON():Ta(a)};Ya=function(a,b){a&128&&Na(b)};
Za=function(a,b,c=Ka){if(null!=a){if(Ca&&a instanceof Uint8Array)return b?a:new Uint8Array(a);if(Array.isArray(a)){const d=_.r(a);if(d&2)return a;if(b&&!(d&32)&&(d&16||0===d))return _.Ga(a,d|18),a;a=Ua(a,Za,d&4?Ka:c,!0,!1);b=_.r(a);b&4&&b&2&&Object.freeze(a);return a}return a.ie===Wa?$a(a):a}};cb=function(a,b,c,d,e,f,g){(a=a.i&&a.i[c])?(d=_.r(a),d&2?d=a:(f=_.ab(a,$a),Ka(d,f),Object.freeze(f),d=f),_.bb(b,c,d,e)):_.t(b,c,Za(d,f,g),e)};
$a=function(a){if(_.r(a.na)&2)return a;a=_.db(a,!0);_.Fa(a.na,18);return a};_.db=function(a,b){const c=a.na;var d=_.Ia([]),e=a.constructor.i;e&&d.push(e);e=a.rb;if(e){d.length=c.length;var f={};d[d.length-1]=f}0!==(_.r(c)&128)&&Na(d);b=b||a.Ib()?Ka:Ja;d=_.Ra(a.constructor,d);a.hd&&(d.hd=a.hd.slice());f=!!(_.r(c)&16);const g=e?c.length-1:c.length;for(let h=0;h<g;h++)cb(a,d,h-a.rc,c[h],!1,f,b);if(e)for(const h in e)cb(a,d,+h,e[h],!0,f,b);return d};
_.eb=function(a){if(!(_.r(a.na)&2))return a;const b=_.db(a,!1);b.s=a;return b};fb=function(a,b){if(Array.isArray(a)){var c=_.r(a),d=1;!b||c&2||(d|=16);(c&d)!==d&&_.Ga(a,c|d)}};gb=function(a,b){return Ta(b)};_.w=function(a,b){return null!=a?!!a:!!b};_.x=function(a,b){void 0==b&&(b="");return null!=a?a:b};_.hb=function(a,b){void 0==b&&(b=0);return null!=a?a:b};
_.jb=function(a,b){let c,d;for(let e=1;e<arguments.length;e++){d=arguments[e];for(c in d)a[c]=d[c];for(let f=0;f<ib.length;f++)c=ib[f],Object.prototype.hasOwnProperty.call(d,c)&&(a[c]=d[c])}};var ob,pb,qb;_.kb=_.kb||{};_.m=this||self;_.lb=function(a,b){a=a.split(".");b=b||_.m;for(var c=0;c<a.length;c++)if(b=b[a[c]],null==b)return null;return b};_.mb=function(a){var b=typeof a;return"object"==b&&null!=a||"function"==b};_.nb="closure_uid_"+(1E9*Math.random()>>>0);ob=function(a,b,c){return a.call.apply(a.bind,arguments)};
pb=function(a,b,c){if(!a)throw Error();if(2<arguments.length){var d=Array.prototype.slice.call(arguments,2);return function(){var e=Array.prototype.slice.call(arguments);Array.prototype.unshift.apply(e,d);return a.apply(b,e)}}return function(){return a.apply(b,arguments)}};_.y=function(a,b,c){Function.prototype.bind&&-1!=Function.prototype.bind.toString().indexOf("native code")?_.y=ob:_.y=pb;return _.y.apply(null,arguments)};
_.z=function(a,b){a=a.split(".");var c=_.m;a[0]in c||"undefined"==typeof c.execScript||c.execScript("var "+a[0]);for(var d;a.length&&(d=a.shift());)a.length||void 0===b?c[d]&&c[d]!==Object.prototype[d]?c=c[d]:c=c[d]={}:c[d]=b};_.B=function(a,b){function c(){}c.prototype=b.prototype;a.V=b.prototype;a.prototype=new c;a.prototype.constructor=a;a.ci=function(d,e,f){for(var g=Array(arguments.length-2),h=2;h<arguments.length;h++)g[h-2]=arguments[h];return b.prototype[e].apply(d,g)}};qb=function(a){return a};
_.rb=function(a){var b=null,c=_.m.trustedTypes;if(!c||!c.createPolicy)return b;try{b=c.createPolicy(a,{createHTML:qb,createScript:qb,createScriptURL:qb})}catch(d){_.m.console&&_.m.console.error(d.message)}return b};_.B(_.ba,Error);_.ba.prototype.name="CustomError";_.sb=function(a){return/^[\s\xa0]*$/.test(a)};_.tb=String.prototype.trim?function(a){return a.trim()}:function(a){return/^[\s\xa0]*([\s\S]*?)[\s\xa0]*$/.exec(a)[1]};var da,ub=_.lb("WIZ_global_data.oxN3nb"),vb=ub&&ub[610401301];da=null!=vb?vb:!1;var wb;wb=_.m.navigator;_.ea=wb?wb.userAgentData||null:null;_.xb=function(a,b){return Array.prototype.indexOf.call(a,b,void 0)};_.yb=function(a,b,c){Array.prototype.forEach.call(a,b,c)};_.ab=function(a,b,c){return Array.prototype.map.call(a,b,c)};_.zb=function(a){_.zb[" "](a);return a};_.zb[" "]=function(){};var Mb,Nb,Sb;_.Ab=_.ia();_.D=_.ja();_.Bb=_.n("Edge");_.Cb=_.Bb||_.D;_.Db=_.n("Gecko")&&!_.ya()&&!(_.n("Trident")||_.n("MSIE"))&&!_.n("Edge");_.Eb=_.ya();_.Fb=_.va();_.Gb=_.wa();_.Hb=_.sa();_.Ib=ta();_.Jb=_.n("iPad");_.Kb=_.n("iPod");_.Lb=_.ua();Mb=function(){var a=_.m.document;return a?a.documentMode:void 0};
a:{var Ob="",Pb=function(){var a=_.ca();if(_.Db)return/rv:([^\);]+)(\)|;)/.exec(a);if(_.Bb)return/Edge\/([\d\.]+)/.exec(a);if(_.D)return/\b(?:MSIE|rv)[: ]([^\);]+)(\)|;)/.exec(a);if(_.Eb)return/WebKit\/(\S+)/.exec(a);if(_.Ab)return/(?:Version)[ \/]?(\S+)/.exec(a)}();Pb&&(Ob=Pb?Pb[1]:"");if(_.D){var Qb=Mb();if(null!=Qb&&Qb>parseFloat(Ob)){Nb=String(Qb);break a}}Nb=Ob}_.Rb=Nb;if(_.m.document&&_.D){var Tb=Mb();Sb=Tb?Tb:parseInt(_.Rb,10)||void 0}else Sb=void 0;_.Ub=Sb;_.Vb=_.ma();_.Wb=ta()||_.n("iPod");_.Xb=_.n("iPad");_.Yb=_.pa();_.Zb=_.na();_.$b=_.oa()&&!_.ua();var ac;ac={};_.bc=null;_.Aa=function(a,b){void 0===b&&(b=0);_.cc();b=ac[b];const c=Array(Math.floor(a.length/3)),d=b[64]||"";let e=0,f=0;for(;e<a.length-2;e+=3){var g=a[e],h=a[e+1],l=a[e+2],q=b[g>>2];g=b[(g&3)<<4|h>>4];h=b[(h&15)<<2|l>>6];l=b[l&63];c[f++]=q+g+h+l}q=0;l=d;switch(a.length-e){case 2:q=a[e+1],l=b[(q&15)<<2]||d;case 1:a=a[e],c[f]=b[a>>2]+b[(a&3)<<4|q>>4]+l+d}return c.join("")};
_.cc=function(){if(!_.bc){_.bc={};for(var a="ABCDEFGHIJKLMNOPQRSTUVWXYZabcdefghijklmnopqrstuvwxyz0123456789".split(""),b=["+/=","+/","-_=","-_.","-_"],c=0;5>c;c++){var d=a.concat(b[c].split(""));ac[c]=d;for(var e=0;e<d.length;e++){var f=d[e];void 0===_.bc[f]&&(_.bc[f]=e)}}}};var Ca;Ca="undefined"!==typeof Uint8Array;_.za=!_.D&&"function"===typeof _.m.btoa;_.dc="undefined"!==typeof TextDecoder;_.ec="undefined"!==typeof TextEncoder;_.Ea=Symbol();var Wa,fc;Wa={};_.gc=Object.freeze(_.Ga([],23));var hc;hc=function(a){const b=a.j+a.rc;return a.rb||(a.rb=a.na[b]={})};_.E=function(a,b,c){return-1===b?null:b>=a.j?a.rb?a.rb[b]:void 0:c&&a.rb&&(c=a.rb[b],null!=c)?c:a.na[b+a.rc]};_.t=function(a,b,c,d){_.Ma(a);return _.ic(a,b,c,d)};_.ic=function(a,b,c,d){a.s&&(a.s=void 0);if(b>=a.j||d)return hc(a)[b]=c,a;a.na[b+a.rc]=c;(c=a.rb)&&b in c&&delete c[b];return a};_.F=function(a,b){a=_.E(a,b);return null==a?a:!!a};
_.jc=function(a,b,c,d){const e=_.E(a,c,d);{let f=!1;null==e||"object"!==typeof e||(f=Array.isArray(e))||e.ie!==Wa?f?(_.Oa(e,_.r(a.na)),b=new b(e)):b=void 0:b=e}b!==e&&null!=b&&_.ic(a,c,b,d);return b};_.G=function(a,b,c,d=!1){b=_.jc(a,b,c,d);if(null==b)return b;if(!(_.r(a.na)&2)){const e=_.eb(b);e!==b&&(b=e,_.ic(a,c,b,d))}return b};_.H=function(a,b,c){_.Ma(a);null==c&&(c=void 0);return _.ic(a,b,c)};
_.bb=function(a,b,c,d){_.Ma(a);var e=null==c?_.gc:_.Ha([]);if(null!=c){var f=!!c.length;for(var g=0;g<c.length;g++){const h=c[g];f=f&&!(_.r(h.na)&2);e[g]=h.na}f=(f?8:0)|1;g=_.r(e);(g&f)!==f&&(Object.isFrozen(e)&&(e=Array.prototype.slice.call(e)),_.Ga(e,g|f));a.i||(a.i={});a.i[b]=c}else a.i&&(a.i[b]=void 0);return _.ic(a,b,e,d)};_.kc=function(a,b,c=0){return _.Pa(_.E(a,b),c)};
_.lc=function(a,b,c=0){const d=_.E(a,b);var e=null==d?d:"number"===typeof d||"NaN"===d||"Infinity"===d||"-Infinity"===d?Number(d):void 0;null!=e&&e!==d&&_.ic(a,b,e);return _.Pa(e,c)};var Qa;_.I=class{constructor(a,b,c){null==a&&(a=Qa);Qa=void 0;var d=this.constructor.i;if(null==a){a=d?[d]:[];var e=!0;_.Ga(a,48)}else{if(!Array.isArray(a))throw Error();if(d&&d!==a[0])throw Error();var f=_.Fa(a,0)|32;e=0!==(16&f);if(128&f)throw Error();_.Ga(a,f)}this.rc=d?0:-1;this.i=void 0;this.na=a;a:{f=this.na.length;d=f-1;if(f&&(f=this.na[d],La(f))){this.rb=f;this.j=d-this.rc;break a}void 0!==b&&-1<b?(this.j=Math.max(b,d+1-this.rc),this.rb=void 0):this.j=Number.MAX_VALUE}if(this.rb&&"g"in this.rb)throw Error("t");
if(c){b=e&&!0;e=this.j;let h;for(d=0;d<c.length;d++)if(f=c[d],f<e){f+=this.rc;var g=a[f];g?fb(g,b):a[f]=_.gc}else h||(h=hc(this)),(g=h[f])?fb(g,b):h[f]=_.gc}}toJSON(){const a=this.na;var b;fc?b=a:b=Ua(a,Xa,Ya,void 0,!1);return b}Fa(){fc=!0;try{return JSON.stringify(this.toJSON(),gb)}finally{fc=!1}}Ib(){return!!(_.r(this.na)&2)}};_.I.prototype.ie=Wa;_.I.prototype.toString=function(){return this.na.toString()};_.mc=Symbol();_.nc=Symbol();_.oc=Symbol();_.pc=Symbol();var qc=class extends _.I{constructor(){super()}};_.rc=class extends _.I{constructor(){super()}rd(a){return _.t(this,3,a)}};_.sc=class extends _.I{constructor(a){super(a)}};var tc=class extends _.I{constructor(a){super(a)}};_.uc=class extends _.I{constructor(a){super(a)}Jc(a){return _.t(this,24,a)}};_.vc=class extends _.I{constructor(a){super(a)}};_.J=function(){this.Ga=this.Ga;this.oa=this.oa};_.J.prototype.Ga=!1;_.J.prototype.isDisposed=function(){return this.Ga};_.J.prototype.ma=function(){this.Ga||(this.Ga=!0,this.N())};_.J.prototype.N=function(){if(this.oa)for(;this.oa.length;)this.oa.shift()()};var wc=class extends _.J{constructor(){var a=window;super();this.o=a;this.i=[];this.j={}}resolve(a){var b=this.o;a=a.split(".");for(var c=a.length,d=0;d<c;++d)if(b[a[d]])b=b[a[d]];else return null;return b instanceof Function?b:null}Uc(){for(var a=this.i.length,b=this.i,c=[],d=0;d<a;++d){var e=b[d].i(),f=this.resolve(e);if(f&&f!=this.j[e])try{b[d].Uc(f)}catch(g){}else c.push(b[d])}this.i=c.concat(b.slice(a))}};var zc=class extends _.J{constructor(){var a=_.yc;super();this.o=a;this.v=this.i=null;this.s=0;this.B={};this.j=!1;a=window.navigator.userAgent;0<=a.indexOf("MSIE")&&0<=a.indexOf("Trident")&&(a=/\b(?:MSIE|rv)[: ]([^\);]+)(\)|;)/.exec(a))&&a[1]&&9>parseFloat(a[1])&&(this.j=!0)}A(a,b){this.i=b;this.v=a;b.preventDefault?b.preventDefault():b.returnValue=!1}};_.Ac=class{constructor(){this.data={}}Fa(a){var b=[],c;for(c in this.data)b.push(encodeURIComponent(c)+"="+encodeURIComponent(String(this.data[c])));return("atyp=i&zx="+(new Date).getTime()+"&"+b.join("&")).substr(0,a)}};var Bc=class extends _.Ac{constructor(a,b){super();var c=_.G(a,tc,8)||new tc;window.google&&window.google.kEI&&(this.data.ei=window.google.kEI);this.data.sei=_.x(_.E(a,10));this.data.ogf=_.x(_.E(c,3));this.data.ogrp=(window.google&&window.google.sn?!/.*hp$/.test(window.google.sn):_.w(_.F(a,7)))?"1":"";this.data.ogv=_.x(_.E(c,6))+"."+_.x(_.E(c,7));this.data.ogd=_.x(_.E(a,21));this.data.ogc=_.x(_.E(a,20));this.data.ogl=_.x(_.E(a,5));b&&(this.data.oggv=b)}};var ib="constructor hasOwnProperty isPrototypeOf propertyIsEnumerable toLocaleString toString valueOf".split(" ");_.Cc=class extends Bc{constructor(a,b,c,d,e){super(a,b);_.jb(this.data,{jexpid:_.x(_.E(a,9)),srcpg:"prop="+_.x(_.E(a,6)),jsr:Math.round(1/d),emsg:c.name+":"+c.message});if(e){e._sn&&(e._sn="og."+e._sn);for(const f in e)this.data[encodeURIComponent(f)]=e[f]}}};var Dc;_.Ec=function(){void 0===Dc&&(Dc=_.rb("ogb-qtm#html"));return Dc};_.Gc=class{constructor(a,b){this.i=b===_.Fc?a:""}toString(){return this.i+""}};_.Gc.prototype.Ab=!0;_.Gc.prototype.hb=function(){return this.i.toString()};_.Ic=function(a){return _.Hc(a).toString()};_.Hc=function(a){return a instanceof _.Gc&&a.constructor===_.Gc?a.i:"type_error:TrustedResourceUrl"};_.Fc={};var Mc,Nc,Qc,Sc,Jc;_.Kc=class{constructor(a,b){this.i=b===Jc?a:""}toString(){return this.i.toString()}};_.Kc.prototype.Ab=!0;_.Kc.prototype.hb=function(){return this.i.toString()};_.Lc=function(a){return a instanceof _.Kc&&a.constructor===_.Kc?a.i:"type_error:SafeUrl"};Mc=/^data:(.*);base64,[a-z0-9+\/]+=*$/i;Nc=/^(?:(?:https?|mailto|ftp):|[^:/?#]*(?:[/?#]|$))/i;
_.Pc=function(a){if(a instanceof _.Kc)return a;a="object"==typeof a&&a.Ab?a.hb():String(a);Nc.test(a)?a=_.Oc(a):(a=String(a).replace(/(%0A|%0D)/g,""),a=a.match(Mc)?_.Oc(a):null);return a};try{new URL("s://g"),Qc=!0}catch(a){Qc=!1}Sc=Qc;
_.Tc=function(a){if(a instanceof _.Kc)return a;a="object"==typeof a&&a.Ab?a.hb():String(a);a:{var b=a;if(Sc){try{var c=new URL(b)}catch(d){b="https:";break a}b=c.protocol}else b:{c=document.createElement("a");try{c.href=b}catch(d){b=void 0;break b}b=c.protocol;b=":"===b||""===b?"https:":b}}"javascript:"===b&&(a="about:invalid#zClosurez");return _.Oc(a)};Jc={};_.Oc=function(a){return new _.Kc(a,Jc)};_.Uc=_.Oc("about:invalid#zClosurez");_.Vc={};_.Wc=class{constructor(a,b){this.i=b===_.Vc?a:"";this.Ab=!0}hb(){return this.i}toString(){return this.i.toString()}};_.Xc=new _.Wc("",_.Vc);_.Yc=RegExp("^[-+,.\"'%_!#/ a-zA-Z0-9\\[\\]]+$");_.Zc=RegExp("\\b(url\\([ \t\n]*)('[ -&(-\\[\\]-~]*'|\"[ !#-\\[\\]-~]*\"|[!#-&*-\\[\\]-~]*)([ \t\n]*\\))","g");
_.$c=RegExp("\\b(calc|cubic-bezier|fit-content|hsl|hsla|linear-gradient|matrix|minmax|radial-gradient|repeat|rgb|rgba|(rotate|scale|translate)(X|Y|Z|3d)?|steps|var)\\([-+*/0-9a-zA-Z.%#\\[\\], ]+\\)","g");var ad;ad={};_.cd=function(a){return a instanceof _.bd&&a.constructor===_.bd?a.i:"type_error:SafeHtml"};_.dd=function(a){const b=_.Ec();a=b?b.createHTML(a):a;return new _.bd(a,ad)};_.bd=class{constructor(a,b){this.i=b===ad?a:"";this.Ab=!0}hb(){return this.i.toString()}toString(){return this.i.toString()}};_.ed=new _.bd(_.m.trustedTypes&&_.m.trustedTypes.emptyHTML||"",ad);_.fd=_.dd("<br>");var hd;_.gd=function(a){let b=!1,c;return function(){b||(c=a(),b=!0);return c}}(function(){var a=document.createElement("div"),b=document.createElement("div");b.appendChild(document.createElement("div"));a.appendChild(b);b=a.firstChild.firstChild;a.innerHTML=_.cd(_.ed);return!b.parentElement});hd=/^[\w+/_-]+[=]{0,2}$/;
_.id=function(a){a=(a||_.m).document;return a.querySelector?(a=a.querySelector('style[nonce],link[rel="stylesheet"][nonce]'))&&(a=a.nonce||a.getAttribute("nonce"))&&hd.test(a)?a:"":""};_.jd=RegExp("^\\s{3,4}at(?: (?:(.*?)\\.)?((?:new )?(?:[a-zA-Z_$][\\w$]*|<anonymous>))(?: \\[as ([a-zA-Z_$][\\w$]*)\\])?)? (?:\\(unknown source\\)|\\(native\\)|\\((?:eval at )?((?:http|https|file)://[^\\s)]+|javascript:.*)\\)|((?:http|https|file)://[^\\s)]+|javascript:.*))$");_.kd=RegExp("^(?:(.*?)\\.)?([a-zA-Z_$][\\w$]*(?:/.?<)?)?(\\(.*\\))?@(?::0|((?:http|https|file)://[^\\s)]+|javascript:.*))$");var ld,od,nd;_.md=function(a){let b;b=window.google&&window.google.logUrl?"":"https://www.google.com";b+="/gen_204?use_corp=on&";b+=a.Fa(2040-b.length);ld(_.Pc(b)||_.Uc)};ld=function(a){var b=new Image,c=nd;b.onerror=b.onload=b.onabort=function(){c in od&&delete od[c]};od[nd++]=b;b.src=_.Lc(a)};od=[];nd=0;_.pd=class extends _.I{constructor(a){super(a)}};_.qd=a=>{var b="wc";if(a.wc&&a.hasOwnProperty(b))return a.wc;b=new a;return a.wc=b};var wd,sd,ud;_.td=function(a,b){var c=_.rd.i();if(a in c.i){if(c.i[a]!=b)throw new sd;}else{c.i[a]=b;if(b=c.j[a])for(let d=0,e=b.length;d<e;d++)b[d].i(c.i,a);delete c.j[a]}};_.vd=function(a,b){if(b in a.i)return a.i[b];throw new ud;};_.rd=class{constructor(){this.i={};this.j={}}static i(){return _.qd(_.rd)}};wd=class extends _.ba{constructor(){super()}};sd=class extends wd{};ud=class extends wd{};var Ad;_.xd=function(a,b){if(a.i){const c=new qc;_.t(c,1,b.message);_.t(c,2,b.stack);_.t(c,3,b.lineNumber);_.t(c,5,1);b=new _.rc;_.H(b,40,c);a.i.log(98,b)}};
Ad=class{constructor(){var a=yd;this.v=zd;this.j=_.hb(_.lc(a,2,.001),.001);this.B=_.w(_.F(a,1))&&Math.random()<this.j;this.A=_.hb(_.kc(a,3,1),1);this.s=0;this.i=this.o=null}log(a,b){_.xd(this,a);try{if(this.B&&this.s<this.A){try{var c=(this.o||_.vd(_.rd.i(),"lm")).s(a,b)}catch(d){c=new _.Cc(this.v,"quantum:gapiBuildLabel",a,this.j,b)}_.md(c);this.s++}}catch(d){}}};var Bd=[1,2,3,4,5,6,9,10,11,13,14,28,29,30,34,35,37,38,39,40,42,43,48,49,50,51,52,53,62,500],Dd=function(a){if(!Cd){Cd={};for(var b=0;b<Bd.length;b++)Cd[Bd[b]]=!0}return!!Cd[a]},Ed=function(a){a=String(a);return a.replace(".","%2E").replace(",","%2C")},Fd=class extends Bc{constructor(a,b,c,d,e){super(a,"quantum:gapiBuildLabel");_.jb(this.data,{oge:c,ogex:_.x(_.E(a,9)),ogp:_.x(_.E(a,6)),ogsr:Math.round(1/(Dd(c)?_.hb(_.lc(b,3,1)):_.hb(_.lc(b,2,1E-4)))),ogus:d});if(e){"ogw"in e&&(this.data.ogw=e.ogw,
delete e.ogw);"ved"in e&&(this.data.ved=e.ved,delete e.ved);a=[];for(var f in e)0!=a.length&&a.push(","),a.push(Ed(f)),a.push("."),a.push(Ed(e[f]));e=a.join("");""!=e&&(this.data.ogad=e)}}},Cd=null;var Gd=class extends _.I{constructor(a){super(a)}};var Kd=class{constructor(){var a=Hd,b=Id,c=Jd;this.j=a;this.i=b;this.s=_.hb(_.lc(a,2,1E-4),1E-4);this.B=_.hb(_.lc(a,3,1),1);b=Math.random();this.o=_.w(_.F(a,1))&&b<this.s;this.v=_.w(_.F(a,1))&&b<this.B;a=0;_.w(_.F(c,1))&&(a|=1);_.w(_.F(c,2))&&(a|=2);_.w(_.F(c,3))&&(a|=4);this.A=a}log(a,b){try{if(Dd(a)?this.v:this.o){var c=new Fd(this.i,this.j,a,this.A,b);_.md(c)}}catch(d){}}};var Md;_.Ld=function(a){if(0<a.o.length){var b=void 0!==a.i,c=void 0!==a.j;if(b||c){b=b?a.s:a.v;c=a.o;a.o=[];try{_.yb(c,b,a)}catch(d){console.error(d)}}}};_.Nd=class{constructor(a){this.i=a;this.j=void 0;this.o=[]}then(a,b,c){this.o.push(new Md(a,b,c));_.Ld(this)}resolve(a){if(void 0!==this.i||void 0!==this.j)throw Error("B");this.i=a;_.Ld(this)}s(a){a.j&&a.j.call(a.i,this.i)}v(a){a.o&&a.o.call(a.i,this.j)}};Md=class{constructor(a,b,c){this.j=a;this.o=b;this.i=c}};_.K=class{constructor(){this.s=new _.Nd;this.i=new _.Nd;this.A=new _.Nd;this.v=new _.Nd;this.B=new _.Nd;this.C=new _.Nd;this.o=new _.Nd;this.j=new _.Nd;this.G=new _.Nd}J(){return this.s}L(){return this.i}M(){return this.A}K(){return this.v}Ga(){return this.B}oa(){return this.C}H(){return this.o}F(){return this.j}static i(){return _.qd(_.K)}};var Sd;_.Pd=function(){return _.G(_.Od,_.uc,1)};_.Qd=function(){return _.G(_.Od,_.vc,5)};Sd=class extends _.I{constructor(){super(Rd)}};var Rd;window.gbar_&&window.gbar_.CONFIG?Rd=window.gbar_.CONFIG[0]||{}:Rd=[];_.Od=new Sd;var yd,zd,Id,Jd,Hd;yd=_.G(_.Od,_.pd,3)||new _.pd;zd=_.Pd()||new _.uc;_.yc=new Ad;Id=_.Pd()||new _.uc;Jd=_.Qd()||new _.vc;Hd=_.G(_.Od,Gd,4)||new Gd;_.Td=new Kd;_.z("gbar_._DumpException",function(a){_.yc?_.yc.log(a):console.error(a)});_.Ud=new zc;_.Td.log(8,{m:"BackCompat"==document.compatMode?"q":"s"});_.z("gbar.A",_.Nd);_.Nd.prototype.aa=_.Nd.prototype.then;_.z("gbar.B",_.K);_.K.prototype.ba=_.K.prototype.L;_.K.prototype.bb=_.K.prototype.M;_.K.prototype.bd=_.K.prototype.Ga;_.K.prototype.bf=_.K.prototype.J;_.K.prototype.bg=_.K.prototype.K;_.K.prototype.bh=_.K.prototype.oa;_.K.prototype.bj=_.K.prototype.H;_.K.prototype.bk=_.K.prototype.F;_.z("gbar.a",_.K.i());var Vd=new wc;_.td("api",Vd);var Wd=_.Qd()||new _.vc;window.__PVT=_.x(_.E(Wd,8));
_.td("eq",_.Ud);
}catch(e){_._DumpException(e)}
try{
_.Xd=class extends _.I{constructor(a){super(a)}};
}catch(e){_._DumpException(e)}
try{
_.Yd=class extends _.I{constructor(a){super(a)}};
}catch(e){_._DumpException(e)}
try{
var Zd=class extends _.I{constructor(){super()}};var $d=class extends _.J{constructor(){super();this.j=[];this.i=[]}o(a,b){this.j.push({features:a,options:b})}init(a,b,c){window.gapi={};var d=window.___jsl={};d.h=_.x(_.E(a,1));null!=_.E(a,12,!1)&&(d.dpo=_.w(_.F(a,12)));d.ms=_.x(_.E(a,2));d.m=_.x(_.E(a,3));d.l=[];_.E(b,1)&&(a=_.E(b,3))&&this.i.push(a);_.E(c,1)&&(c=_.E(c,2))&&this.i.push(c);_.z("gapi.load",(0,_.y)(this.o,this));return this}};var ae=_.G(_.Od,_.Xd,14)||new _.Xd,be=_.G(_.Od,_.Yd,9)||new _.Yd,ce=new Zd,de=new $d;de.init(ae,be,ce);_.td("gs",de);
}catch(e){_._DumpException(e)}
})(this.gbar_);
// Google Inc.
</script><title>LAB03</title><script nonce="">var AF_initDataKeys = []; var AF_dataServiceRequests = {}; var AF_initDataChunkQueue = []; var AF_initDataCallback; var AF_initDataInitializeCallback; if (AF_initDataInitializeCallback) {AF_initDataInitializeCallback(AF_initDataKeys, AF_initDataChunkQueue, AF_dataServiceRequests);}if (!AF_initDataCallback) {AF_initDataCallback = function(chunk) {AF_initDataChunkQueue.push(chunk);};}</script><script async="" type="text/javascript" charset="UTF-8" src="dec2_to_4_files/rs=AA2YrTvkbJWV1adPbuzYq0DsgPYnetf7Bg" nonce=""></script><link type="text/css" rel="stylesheet" href="dec2_to_4_files/rs=AA2YrTvmtKM57xcbKdJeX3djH0NMhQr_Nw.css" nonce=""><style nonce="" type="text/css" data-late-css="">.hD8oBb.hD8oBb,.hD8oBb .T4LgNb{height:100%}.hD8oBb .kFwPee{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;height:100%;overflow:hidden}@media (max-width:30rem){.hD8oBb .kFwPee{height:auto}}.C7gDne{display:-moz-box;display:flex;-moz-box-flex:1;flex:1 1 auto;-moz-box-pack:center;justify-content:center;overflow:hidden}@media (max-width:30rem){.C7gDne{display:block}}.mI0dk{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;overflow:hidden}.SbtHLc{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;padding:1rem 1rem 0}@media not all and (max-width:61.25rem){.i3Utwc{-moz-box-flex:0;flex:0 1 33.3333333333%}}@media (max-width:61.25rem){.SbtHLc{-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.F9zdgb{align-self:flex-start;margin-bottom:1rem}}.SqncUb{display:-moz-box;display:flex;-moz-box-pack:center;justify-content:center;padding:.75rem;margin:-.75rem}.CFcF2d{display:inline-block;text-align:center;margin:0 1rem;min-width:9.5rem}.V203cd{border-radius:px-to-rem(4);display:-moz-box;display:flex;-moz-box-flex:1;flex:1 1 auto;overflow:auto;margin:1rem;margin-bottom:1.5rem;max-width:calc(100vw - 2.125rem)}.gYzugb{visibility:hidden}.RIDjNe{border-right:.0625rem solid rgb(218,220,224);-moz-box-sizing:border-box;box-sizing:border-box;display:-moz-box;display:flex;-moz-box-flex:0;flex:0 0 10.5357142857rem;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;font-weight:500;overflow:hidden;width:10.5357142857rem}.RIDjNe:last-child{border-right:0}.yAAeVc{overflow-y:auto}.dYwBL{border-radius:.125rem;display:block;margin:.25rem;padding:.5rem;text-decoration:none;word-wrap:break-word}.MjKYZc{color:#fff;font-weight:500}.THta6c{color:#fff;font-weight:400}.Eajscb{display:-moz-box;display:flex;-moz-box-pack:center;justify-content:center;padding-bottom:1.5rem}.Eajscb .vT1Gyc{border-radius:100%;height:2.875rem;line-height:2.875rem;margin-top:-.5rem;text-align:center;width:2.875rem}.Eajscb .vT1Gyc.pCcXPe{color:#70757a}.Eajscb .vT1Gyc.F262Ye{background-color:rgb(26,115,232);color:#fff}.Eajscb .vT1Gyc.N4XV7d{color:rgb(60,64,67)}.Eajscb .nGZbac,.Eajscb .nGZbac.pCcXPe,.Eajscb .nGZbac.N4XV7d{color:#70757a;line-height:2rem;margin-left:0;margin-top:.5rem;text-align:center}.Eajscb .nGZbac.F262Ye{color:rgb(26,115,232)}.F9zdgb{line-height:1;width:100%}.s8jIAb{color:rgba(0,0,0,.549);margin-right:1rem;text-align:right}.WD0wFe{display:block}@media (max-width:30rem){.V203cd{-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.RIDjNe{border-right:none;display:-moz-box;display:flex;margin-bottom:.5rem;padding:0 1rem 0 1.5rem;width:unset}.yAAeVc{display:-moz-box;display:flex;-moz-box-flex:1;flex:1 1 auto;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.dYwBL{margin-left:0;margin-right:.5rem}.Eajscb{flex-basis:2.5rem;flex-shrink:0;-moz-box-pack:start;justify-content:flex-start;padding-bottom:0;padding-right:.5rem}.Eajscb .vT1Gyc{font-size:1.5rem}.Eajscb .vT1Gyc.F262Ye{background-color:#fff;color:rgb(26,115,232)}.Eajscb .vT1Gyc,.Eajscb .nGZbac,.Eajscb .nGZbac.pCcXPe,.Eajscb .nGZbac.N4XV7d{margin-left:0;text-align:left}}.t4j4Wb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.a3p7rb{width:21.25rem}.CJXzee{flex-shrink:0;margin:0 -1.5rem -1.5rem -1.5rem;overflow:hidden;padding:3.375rem 3.375rem 0.5rem 1.5rem;width:10.125rem}.aJiAfb{font-style:italic}.CJXzee .fXuRkd{align-items:stretch}.CJXzee a{display:block;box-flex:1;flex-grow:1;line-height:3rem;padding-right:1.5rem;position:relative;text-decoration:none}.zFfAHb{padding-left:0.75rem}.CJXzee a:active,.CJXzee a:focus,.CJXzee a:hover{color:rgba(0,0,0,.87);text-decoration:none}.CJXzee a:active .ULzZ3{animation:hrRippleTransform .2s cubic-bezier(0,0,0.2,1) forwards;opacity:.08}.fXuRkd:hover,.zFfAHb:focus{-moz-border-radius:0.5rem;border-radius:0.5rem}.CJXzee a.rUnD6d{font-weight:500;color:inherit;text-decoration:none}.cizThc,.BYOike{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:500}.ByX3Cc{left:1.5rem;position:sticky;width:17.5rem}.DPt8E{min-width:17.5rem}.Tq5Atc{margin:12.5rem auto 0;text-align:center}.nViTIe{height:8.75rem}.UGLIMe{margin:2rem auto .25rem;width:20rem}.w3wv2b{margin-top:1rem}.whsmod{margin-bottom:11.25rem;margin-top:-12.5rem;text-align:left}@media (max-width:40rem){.Tq5Atc{margin-top:6.25rem}.whsmod{margin-bottom:5rem;margin-top:-6.25rem}}.EwF03c{background-color:#fff;border-bottom:.0625rem solid rgb(218,220,224);-moz-box-sizing:border-box;box-sizing:border-box;flex-wrap:nowrap;-moz-box-pack:justify;justify-content:space-between;left:0;padding:.5rem 1.5rem;position:sticky;top:4.0625rem;width:100vw;z-index:5}@media (max-width:65.125rem){.EwF03c{top:8.0625rem}}.rGxdsf{margin-right:-0.875rem}.CmLZs{align-items:flex-start;box-flex:0;flex-grow:0;flex-shrink:0}.a0BN6e.a0BN6e{display:block}.kcAzD:focus:before{border:solid 0.0625rem #9e9e9e;bottom:0;content:" ";left:0;position:absolute;right:0;top:0}.k91PN{table-layout:fixed}.n9BHJf table{border-collapse:collapse;border-spacing:0;height:1px;overflow:hidden;position:relative;table-layout:fixed}.n9BHJf th{height:100%;padding:0}.n9BHJf td{height:100%;padding:0;position:relative}.xZgFJd{width:100%}.vvqDLc{border-bottom:0.0625rem solid #e0e0e0;box-sizing:border-box;height:100%}.go6aXd,.fum4Tb,tbody .vvqDLc{background:#fff}.go6aXd.xAKnLc,.fum4Tb.xAKnLc,tbody .vvqDLc.xAKnLc{background:#f8f9fa}.fHar6b,.RUkyfb,thead .vvqDLc{background:#fff}.n9BHJf th{position:relative;z-index:2}.n9BHJf thead th:first-child{z-index:3}.n9BHJf tbody th:first-child{z-index:1}.n9BHJf th{font-weight:inherit}.fHar6b,.RUkyfb,.go6aXd{box-sizing:border-box;border-bottom:0.0625rem solid #e0e0e0;border-right:0.0625rem solid #e0e0e0;height:100%}.fum4Tb{box-sizing:border-box;border-bottom:0.0625rem solid #e0e0e0;border-right:0.0625rem solid #e0e0e0}.CAdcCb .fHar6b:after{height:110vh;-moz-box-shadow:0px 5px 8px 0px rgba(0,0,0,.14),0px 1px 14px 0px rgba(0,0,0,.12),0px 3px 5px -1px rgba(0,0,0,.2);box-shadow:0px 5px 8px 0px rgba(0,0,0,.14),0px 1px 14px 0px rgba(0,0,0,.12),0px 3px 5px -1px rgba(0,0,0,.2);content:"";pointer-events:none;position:absolute;right:0;top:-5vh;width:100vw;z-index:-1}.RUkyfb{padding:0.75rem 1rem;text-align:left;vertical-align:top}.YV4zId{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.RUkyfb,.fum4Tb{width:8.0625rem}.uzT1Pd{line-height:1.25rem;height:2.5rem;overflow:hidden;text-overflow:ellipsis;word-break:break-word;display:block;display:-webkit-box}.N8tCm .uzT1Pd{overflow:visible}.Pbki4b.O0HS9e:before{border-top:0.0625rem solid #e0e0e0;content:"";display:block}.Pbki4b:before,.YV4zId{padding-bottom:0.25rem}.tpSpse{color:rgba(0,0,0,.549)}.fHar6b{align-items:flex-end;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.N8HYTb{padding-left:3.5rem;padding-right:1.5rem;min-width:11.875rem}.go6aXd{justify-content:space-between}.XnWe0e{padding:0 0.5rem 0 1.5rem}.OnK3U{line-height:2rem;padding-bottom:0.5rem;text-align:left;width:7.0625rem}.tpSpse{text-align:left;width:7.0625rem}.HSanvb{align-self:center;height:2rem;margin-right:1rem;width:2rem}.NhkgIc{font-size:1.5rem;margin-right:1rem;padding:0.25rem}.fum4Tb{height:4rem}.Ws95y{padding:0 1rem}.Y0qupd .n9BHJf .PDpaTd{cursor:pointer}.N8tCm{display:none}.n9BHJf.JpY6Fd .N8tCm{display:table-cell}.pKbqce{cursor:default}.pKbqce:focus:before,.xAKnLc:focus:before{border:solid 0.0625rem #9e9e9e;bottom:0;content:" ";left:0;position:absolute;right:0;top:0}.C31U3e{-moz-box-flex:1 1;flex:1 1;min-width:0}.zIKt9b .RLRLxb .JRtysb{color:transparent}.RUkyfb:hover .RLRLxb .JRtysb,.RUkyfb:focus .RLRLxb .JRtysb,.RLRLxb .JRtysb.iWO5td,.RLRLxb .JRtysb:focus{color:#444}.WAGvmf{max-width:11.875rem}.LCRwqc{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;justify-content:center;width:3.375rem}.L2dBdc{width:100%}.i4mSrb{padding-bottom:0.25rem;width:100%}.CqN3rc{white-space:nowrap}.LCRwqc .MQL3Ob{flex-shrink:0}.w1T5Ae{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;width:100%}.xJVELb{font-style:italic}.S2hMh{margin:0 0.5rem}.LCRwqc .A37UZe{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;padding-left:0}.LCRwqc .oJeWuf{height:auto;width:100%}.LCRwqc .aXBtI{align-items:center;top:0}.LCRwqc .zHQkBf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:0.875rem;font-weight:500;line-height:1.25rem;text-align:right;width:100%}.i4mSrb .snByac{font-size:0.8125rem;line-height:1.25rem;right:0;top:0}.LCRwqc .rFrNMe.u3bW4e .ndJi5d{display:none}.Jqkezb{margin-bottom:0.5rem}.Ek8Cib{height:3.5rem}.xiFNYc{margin-top:0.5rem}.uPXIg .tkmmwb{margin-right:0.5rem;align-self:center}.wmjvHb{text-align:right}.PDpaTd{position:relative}.hDVLxe{overflow:hidden;box-flex:1;flex-grow:1;transition:opacity 0.28s cubic-bezier(0.4,0,0.2,1)}.rRimpd{box-flex:1;flex-grow:1;transition:opacity 0.28s cubic-bezier(0.4,0,0.2,1)}.hDVLxe{opacity:0}.rRimpd{position:absolute}.i5aS4e .rRimpd{opacity:0}.hDVLxe .DPvwYc{display:block}.i5aS4e .hDVLxe{opacity:1}.PDpaTd{height:100%}.gRisWe{height:100%;overflow:hidden;padding:0 1rem;text-overflow:ellipsis}.WLsCn{cursor:text}.oFj0xc{cursor:default}.cL8LOd{border-bottom:0.0625rem solid rgba(0,0,0,.87);display:inline-block;line-height:1;vertical-align:top;width:1.25rem}.EhRlC .cL8LOd{border-bottom-color:#1e8e3e}.lYU7F .cL8LOd{border-bottom-color:#c5221f}.PDpaTd .neggzd.asQXV{color:transparent}.PDpaTd:hover .foVBo,.PDpaTd.Rt1Pjf .foVBo{font-size:0.0625rem;height:0.0625rem;line-height:1;opacity:.001;overflow:hidden;position:absolute;width:0.0625rem}.PDpaTd:not(:hover):not(.Rt1Pjf) .NhG04b{display:none}.PDpaTd.Rt1Pjf:before{border:solid 0.0625rem #9e9e9e;bottom:0;content:" ";left:0;position:absolute;right:0;top:0}.UNDeAc{margin-left:-1rem;margin-right:-0.875rem}.w3SmKe{display:block;font-style:italic}a.qBkhTe{text-decoration:none}.qyDPcd{flex-direction:row-reverse;width:100%}.zCN7Sd{margin-right:1rem}.r9IELc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-shrink:0}.dKqQzd .XEeo8c{border-bottom-right-radius:0;border-top-right-radius:0}.O0rVrc{border-bottom-left-radius:0;border-top-left-radius:0;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-left:-0.0625rem;min-width:2.125rem}.O0rVrc.iWO5td{border-left:1px solid transparent}.O0rVrc .snByac{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.O0rVrc .Fxmcue,.O0rVrc.iWO5td .Fxmcue{padding:0 0.25rem}.O0rVrc .MbhUzd{left:50%!important;top:50%!important}.FiqQZc{transform:scaleX(-1)}.ccG3qf{animation:exportButtonIconSpin 2s linear infinite}@keyframes exportButtonIconSpin{0%{transform:scaleX(-1) rotate(360deg)}to{transform:scaleX(-1) rotate(0deg)}}.wvERWc{color:#b31412;margin-right:0.5rem}.NKcaye{margin-left:1rem}.RGgeHf{height:auto;margin-top:0.625rem;overflow:visible}.RGgeHf .oJeWuf{height:auto;white-space:normal}.RGgeHf .jO7h3c{align-self:center}.ZtITRc{margin:-4px -12px}.XNIQbd{border-collapse:collapse;width:100%}.gQZxn{border:0.0625rem solid #e0e0e0;padding:0.5rem}.e9Ekud{color:rgba(0,0,0,.549);padding:1.5rem}.KTpuI{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.Hn01xe,.Qv6pvf{margin-top:1rem}.k6bWY{display:inline-block;vertical-align:middle}.Era2ub{justify-content:space-between;margin-bottom:0.25rem;padding-left:1rem}.Oo2pXc{position:relative}.Oo2pXc .gQZxn{border-width:0}.ycbm1d{border-top:0.0625rem solid #e0e0e0;height:3.75rem}.ycbm1d:first-child{border-top:0}.p4BDke .ycbm1d:first-child{border-top:0.0625rem solid #e0e0e0}.FvI3qc .d64Ge{padding:0.5rem 1.5rem;text-align:right}.d64Ge .oxacD{display:inline-block}.YG03qb{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:flex-end}.YG03qb .TpQm9d{color:inherit}.zuJ3be{vertical-align:bottom}.T0H2Fb{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.ZDe7q{-moz-box-flex:0 0 2.5rem;flex:0 0 2.5rem;padding:0 0.5rem;text-align:center}.sCv5Q{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;margin-left:0.5rem;max-width:30rem}.ch1JNd .ZDe7q,.ch1JNd .sCv5Q{opacity:0.54}.pXwmie{margin-left:0.5rem}.DKlFId tr{height:3.125rem}.DKlFId td{text-align:center}.G4LVac{padding:0.5rem 1.5rem 0 0;margin-bottom:-0.25rem}@media (max-width:40em){.sCv5Q{max-width:11.25rem}.G4LVac{padding-right:1rem;margin-bottom:0.25rem}.FvI3qc .d64Ge{padding-right:1rem}}.vgNHOd{margin:0.5rem 1rem}.ZbZ7Ne{margin-bottom:0.5rem}.ZbZ7Ne:first-child{margin-top:0.5rem}.TXziZ{padding-left:0.5rem}.I5jije{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.tggdAd{margin:0}.PlhAnc{display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;vertical-align:middle}.HTxhwc .XNIQbd{table-layout:fixed}.HTxhwc .gQZxn{border-width:0}.XxEA4d{box-shadow:0 .0625rem .125rem rgba(0,0,0,.12),0 0 .0625rem rgba(0,0,0,.12)}.d6CWTd{border-top:.0625rem solid rgb(218,220,224);height:3.75rem}.hhj3ub .d6CWTd:not(.Zolage),.hhj3ub .d6CWTd:not(.Zolage) .YHVwkf{cursor:pointer}.XxEA4d{box-shadow:none}.d6CWTd td:first-child{border-top-left-radius:.5rem;border-bottom-left-radius:.5rem}.d6CWTd td:last-child{border-top-right-radius:.5rem;border-bottom-right-radius:.5rem}.hhj3ub .d6CWTd:not(.Zolage):hover,.hhj3ub .d6CWTd:not(.Zolage):hover+.d6CWTd{border-color:transparent}.d6CWTd:first-child{border-top:0}.Zolage .zrBYj,.Zolage .PNAi9e,.Zolage .y4ihN{opacity:.54}.qRU9Ec .DnNMBb{display:none}.wIfvCd{text-align:left}.tjHubc{padding-top:.875rem;vertical-align:top}.tjHubc.Mlpuof{padding-top:1.125rem}.paYY4e{cursor:default;padding:0 0 1rem 0}.NO7Twd{margin-left:.75rem}.iMLbRe,.mdcmqc{font-weight:normal;padding:0 .5rem}.iMLbRe{padding:0 0 0 .5rem}.mdcmqc{padding:0}.mdcmqc .oJeWuf{color:rgba(0,0,0,.549)}.QCzpmc{-moz-box-pack:end;justify-content:flex-end;width:100%}.g2DEGd{padding:0 .5rem;vertical-align:middle}.zrBYj{display:inline-block;-moz-box-flex:0;flex:0 0 3.5rem;padding:0;text-align:center;width:3.5rem}.ofWlVd{margin-left:.5rem}.njrcAb{width:5rem}.PNAi9e{-moz-box-flex:0;flex:0 0 2.5rem;text-align:center;width:2.5rem}.L2QUBc{height:2rem;width:2rem}.WMtsmc{margin:-1rem;overflow:hidden;padding:1rem}.KnNDJe{padding:.75rem 0}.KnNDJe .ofWlVd{display:block}.lkqKH .ofWlVd{display:none}.PeKgHf{padding-right:1rem;text-align:right}.PeKgHf .mUbCce{vertical-align:middle}.DikUaf{padding-right:1.5rem;text-align:right}@media (max-width:40rem){.DikUaf{padding-right:1rem}}.VHfpDb{margin-left:1.5rem}.u5Sz3b{color:rgba(0,0,0,.549);font-weight:500;margin-right:.5rem;text-transform:uppercase}.FSRX6{color:rgba(0,0,0,.549);font-size:.8125rem;font-weight:500;line-height:1rem;margin-left:.5rem;max-width:100%}@media not all and (max-width:40rem){.FSRX6{width:40%}}.YHVwkf{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-flex:1;flex-grow:1;overflow:hidden;height:3.25rem;margin:-.625rem;margin-right:0;padding-left:.625rem}.Mlpuof{padding:.5rem 1.5rem;text-align:right;width:4rem}@media (max-width:40rem){.Mlpuof{padding:0 .5rem 0 0}}.HTxhwc th.Mlpuof{padding:0 1.5rem 1.5rem 1.5rem}.Mlpuof .oxacD{display:inline-block}.Mlpuof .TpQm9d{color:inherit}.WbqQDb{display:-moz-box;display:flex;-moz-box-flex:1;flex-grow:1;flex-wrap:wrap;margin-right:.5rem;overflow:hidden}.KwqU3e{margin-left:.5rem;overflow:hidden;padding:0}@media not all and (max-width:40rem){.iCr7o{width:auto}}@media (max-width:40rem){.d6CWTd td{border-radius:.5rem}.y4ihN{max-width:8.75rem}.iFGZdc{width:100%}.L7xZwf{width:0}.zrBYj{flex-basis:2rem;width:2rem}.xukHhe{display:-moz-box;display:flex;margin-left:4rem;margin-right:1rem}}.MwhM8b{margin-bottom:1rem;padding-left:1rem}.anlSm{display:-moz-box;display:flex;-moz-box-flex:1;flex-grow:1;flex-wrap:wrap;-moz-box-align:baseline;align-items:baseline}.lIPLbd{padding:.5rem 1.5rem 0 0;margin-bottom:-.25rem}.jg22B{padding-right:1.5rem}@media (max-width:40rem){.lIPLbd{padding-right:1rem;margin-bottom:.25rem}.jg22B{padding-right:1rem}}.CPYzFb.MAdsVd .MwhM8b,.hhj3ub.MAdsVd .jg22B{display:none}.t5QO8d{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.ueXqmb{height:8.4375rem;margin-top:6.25rem}@media (max-width:40em){.ueXqmb{margin-top:1.875rem}}.LY7xXe{margin:2rem 0 0.25rem 0}.m3igGd{display:block}.ScTWW{margin-top:-20px}.A5u8bf{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;margin-top:4rem}.FEIuWc{height:10rem}.uSlvFd{margin-top:1.5rem;text-align:center;width:16.875rem}.xBIR3c{margin-bottom:1rem}.xBIR3c:not(.Uy7ePe){cursor:pointer}.xBIR3c.Uy7ePe.YRdPTb .hYsg7c:not(.N2RpBe){visibility:hidden}.xBIR3c .snByac{letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:0.75rem;font-weight:400;line-height:1rem;color:#5f6368}.jZrWoe{margin-bottom:1rem}.jZrWoe:not(:empty){word-wrap:break-word}.tHymfc{padding-bottom:1rem}.uQ3ESd{background-color:white}.NoUlnb,.TaY5Vd{overflow-y:auto}.NoUlnb{max-height:45rem}.TaY5Vd.TaY5Vd{padding-bottom:0}.NoUlnb .e3aEUd{padding:0 1.5rem}.TaY5Vd .e3aEUd{margin-bottom:1rem}.TaY5Vd .e3aEUd.TL3Rwd{margin-bottom:0.75rem;padding-bottom:0.25rem}.NoUlnb .wBxtkd{margin-bottom:1.5rem;padding-top:1.5rem;padding-bottom:0.5rem}.uQ3ESd .aHTZpf{padding-top:0}.NoUlnb .SObBRb{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;height:6.75rem;justify-content:center;margin:0}.CwBXrb{overflow:hidden}.TaY5Vd .CwBXrb{margin-bottom:0}.VDj5V{border-top:0.0625rem solid #e0e0e0;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;padding:0.5rem 1.5rem}.P02DYb{border-top:0.0625rem solid #e0e0e0;height:3.75rem;padding:0 1rem}.TaY5Vd .aHTZpf,.TaY5Vd .VvAAB{margin:0 -1.5rem}.NoUlnb .VvAAB{padding-bottom:1rem}@media (max-width:40em){.NoUlnb{max-height:inherit}}.HG7HUc{padding:0 1.5rem}.aSG3qe{-moz-box-flex:0 0 52%;flex:0 0 52%;overflow:hidden}.Ag63Pe,.cpvBkb,.xw0Qof{-moz-box-flex:0 0 calc(16% - 0.5rem);flex:0 0 calc(16% - 0.5rem)}.Ag63Pe,.cpvBkb{margin-left:0.5rem}.XREa9d{-moz-box-flex:0 0 60%;flex:0 0 60%;overflow:hidden}.edG9I{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.LxYeeb,.Sk7ko{-moz-box-flex:0 1 auto;flex:0 1 auto;max-width:50%}.Sk7ko:not(:empty):before{content:"\002022";display:inline-block;margin:0 0.25rem}@media (max-width:40em){.xw0Qof{-moz-box-flex:0 0 calc(40% - 0.5rem);flex:0 0 calc(40% - 0.5rem)}}.xw0Qof{text-align:right}@media (max-width:30em){.HG7HUc{padding:0 0.5rem}}.MZx95d:not(:empty){margin-left:0.75rem}.aP1Rbb{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.sr2FGb{box-flex:1;flex-grow:1;margin-right:0.5rem 1rem 0 1rem;padding:0 0 0 1.5rem}.rVhh3b{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;margin-bottom:1.5rem}@media (max-width:40em){.n0bz1e{margin:0;margin-top:1.5rem;width:100%}}@media (max-width:30em){.n0bz1e{margin:0}}.XU2Svc{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding-bottom:4rem;padding-top:4rem}.U1RWTe .f0kHoc{padding-top:4rem}.i1wJG{padding-top:0}.ts0Nhe{align-items:center;box-sizing:border-box;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.i1wJG.uO32ac{height:auto}.xeNpM{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;width:100%}.YEvYV{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-top:1rem;width:100%}.DIZjNc{-moz-border-radius:50%;border-radius:50%;flex-shrink:0;height:4.6875rem;width:4.6875rem}.qp1Eye{overflow:hidden}.vNFzIf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:2.25rem;font-weight:400;line-height:2.75rem;cursor:pointer}.UJPoPd{display:none}@media not all and (max-width:40em){.DIZjNc{margin-right:1.5rem}}@media (max-width:40em){.ts0Nhe{flex-direction:column}.qp1Eye{align-self:stretch}}.F3Fywc{margin-right:1rem}.yPbwG{align-items:center;-moz-border-radius:0;border-radius:0;margin-bottom:1.5rem;max-width:100%}.sPtISb{-moz-border-radius:0;border-radius:0;padding:0.5rem 1rem;padding-right:0.5rem;text-align:left;width:100%}.sPtISb.RDPZE .snByac{opacity:.54}.sPtISb .snByac{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;width:100%}.sPtISb .Fxmcue{padding:0}.Pxfnyf.Pxfnyf{align-self:center;margin-right:1rem}.xN4Z8e{overflow:hidden}.ECOutf{box-sizing:border-box;padding:1.5rem;width:100%}.WdYux{color:#7f7f7f;font-size:0.875rem;margin-bottom:0.5rem}.cY2sGe{margin-top:0.5rem}.OIh3D{flex-flow:row wrap}.tWKJ2{margin-top:1rem}.RnC9kd{margin:0 0 0.5rem 1rem}.Ti8cTc{max-width:100%;width:29rem}.JB501c{display:table}.KhAuve{display:table-row}.wPGir{color:#7f7f7f;display:table-cell}.utxoK,.rsDI7e,.VvshNc{display:table-cell;overflow:hidden;white-space:normal;word-break:break-word}.utxoK,.rsDI7e{font-weight:500;padding-left:16px}.PpfbXd{padding-top:0.5rem}.VvshNc{vertical-align:top}.VvshNc .LMgvRb .oJeWuf{max-width:9.75rem}.VvshNc .OA0qNb .oJeWuf{text-overflow:ellipsis;overflow:hidden;white-space:nowrap;display:block;max-width:22.5rem}@media (max-width:40em){.VvshNc .LMgvRb .oJeWuf{font-size:0.875rem}}.KojGNd{margin:1rem 0}.RwArwf{display:block;max-width:100%;overflow-y:auto}.RwArwf>.oJeWuf{overflow-y:visible}.aahm2d{padding-bottom:0.5rem}.aahm2d:not(:last-child){border-bottom:0.0625rem solid #e0e0e0;margin-bottom:1.5rem}.KbCMnb{margin:0.5rem 0 0.5rem 3.5rem}.hDBexb{overflow:hidden}.XSCXFb{margin:1rem 0;max-width:100%;width:20rem}.ylfEac{border-bottom:0.0625rem solid #e0e0e0}.nd18Yd{overflow:visible}.VXX6Hf{padding:1.5rem 1.5rem 0}.SCzU2e{margin-bottom:1.5rem}.ripncc{margin-bottom:0.5rem}@media (max-width:48.75em){.QxHFHb{margin:0 1rem}.SCzU2e{margin-bottom:0.5rem}}.VeJ8me.VeJ8me.VeJ8me{max-width:24rem}.JRosVd{color:white}.fCTDtb,.fCTDtb:hover{opacity:.15}.eaBpBc{animation:hrCourseDriveIconFadeIn .5s}.xp2dJ .eaBpBc{animation:none}@keyframes hrCourseDriveIconFadeIn{0%{opacity:.15}to{opacity:0.54}}.gHz6xd{background-clip:padding-box;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;height:18.375rem;margin-bottom:1.5rem;margin-right:1.5rem;overflow:hidden;position:relative;text-align:left;width:18.75rem}.gHz6xd.KQjUpc:hover{box-shadow:0 8px 10px 1px rgba(0,0,0,.14),0 3px 14px 2px rgba(0,0,0,.12),0 5px 5px -3px rgba(0,0,0,.2)}.gHz6xd.xp2dJ{box-shadow:0 8px 10px 1px rgba(0,0,0,.14),0 3px 14px 2px rgba(0,0,0,.12),0 5px 5px -3px rgba(0,0,0,.2);cursor:move;opacity:.9}.TisIWb .kKn9Nc,.TisIWb .kKn9Nc:hover{background-color:transparent;border-color:transparent;box-shadow:none;position:relative;visibility:visible}.TisIWb .kKn9Nc *{visibility:hidden}.TisIWb .kKn9Nc:before{background-color:rgb(241,243,244);bottom:0;content:"";left:0;position:absolute;right:0;top:0;z-index:0}@media (max-width:40rem){.TisIWb .TQYOZc,.TisIWb .SZ0kZe,.TisIWb .F2CcI,.xp2dJ .TQYOZc,.xp2dJ .SZ0kZe,.xp2dJ .F2CcI{display:none}.TisIWb .gHz6xd,.gHz6xd.xp2dJ{border:none;height:auto}}.gHz6xd.rZXyy:not(.kKn9Nc):not(.u0dx8e):hover{border:none;margin:.0625rem 1.5625rem 1.5625rem .0625rem}.OoQyKf{opacity:.5}.Tc9hUd{position:relative}.OjOEXb,.ZizeYd,.O7utsb,.ZmqAt{height:100%;left:0;position:absolute;top:0;width:100%}.OjOEXb{background-repeat:no-repeat;background-size:cover}html[dir=rtl] .OjOEXb.Gf8MK{transform:scaleX(-1)}.ZizeYd{background-color:#999;opacity:.8}.ZizeYd{opacity:.7}.ZizeYd,.O7utsb{background-color:rgb(32,33,36)}.R4EiSb{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-pack:justify;justify-content:space-between;height:4.5rem;padding:1rem 1rem .75rem;position:relative}.lJv9ke{-moz-box-flex:0;flex:0 0 4.6875rem}.prWPdf{display:-moz-box;display:flex;color:white}.prWPdf,.jJIbcc{position:relative}.eDfb1d{display:block;margin:0 -.25rem;padding:0 .25rem}.PNzAWd{border-radius:50%;float:right;height:4.6875rem;position:relative;margin-top:-3.09375rem;width:4.6875rem}.TQYOZc{-moz-box-flex:1;flex-grow:1;min-height:0;padding:1rem;padding-top:.75rem}.TQYOZc .sdDCme{display:none}.F2CcI,.SZ0kZe{display:-moz-box;display:flex;flex-shrink:0;-moz-box-pack:end;justify-content:flex-end}.F2CcI{padding:1rem}.F2CcI{padding:.5rem 1rem}.SZ0kZe{border-top:.0625rem solid rgb(218,220,224);line-height:0;padding:.25rem}.BnYgFe{background-image:-webkit-repeating-linear-gradient(-135deg,transparent,transparent .5625rem,rgba(255,255,255,.3) .5625rem,rgba(255,255,255,.3) .625rem);background-image:repeating-linear-gradient(-135deg,transparent,transparent .5625rem,rgba(255,255,255,.3) .5625rem,rgba(255,255,255,.3) .625rem);background-size:.8838834765rem .8838834765rem;bottom:-50%;left:-50%;pointer-events:none;position:absolute;right:-50%;top:-50%;transform:rotateZ(15deg)}a.kj3hr:hover,a.kj3hr:focus,a.kj3hr:visited{color:#fff}a.kj3hr:focus{background-color:rgba(255,255,255,.25);border-radius:.125rem}.JwPp0e{display:-moz-box;display:flex;flex-wrap:wrap;padding-left:1.5rem;padding-top:1.5rem}.VMO3ed{margin-left:1.5rem;margin-top:1.5rem;width:18.75rem}.VMO3ed .KC1dQ{border-color:transparent}.zOIsg{background-color:rgb(248,249,250);height:100%;width:100%;padding:1rem}.Udkveb{display:-moz-box;display:flex}.giBm9d{height:2.5rem;width:2.5rem;border-radius:50%;background-color:rgb(232,234,237)}.oTdC6b{margin:.5rem}.raAzUc{margin:auto .5rem}.VSG5Ac{margin:.5rem;margin-left:auto}.eut1lf{margin-top:1rem;position:relative}.VfPpkd-WsjYwc{border-radius:4px;border-radius:var(--mdc-shape-medium,4px);background-color:#fff;background-color:var(--mdc-theme-surface,#fff);position:relative;box-shadow:0 2px 1px -1px rgba(0,0,0,.2),0 1px 1px 0 rgba(0,0,0,.14),0 1px 3px 0 rgba(0,0,0,.12)}.VfPpkd-WsjYwc .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-WsjYwc::after{border-radius:4px;border-radius:var(--mdc-shape-medium,4px)}.VfPpkd-WsjYwc-OWXEXe-INsAgc{box-shadow:0 0 0 0 rgba(0,0,0,.2),0 0 0 0 rgba(0,0,0,.14),0 0 0 0 rgba(0,0,0,.12);border-width:1px;border-style:solid;border-color:#e0e0e0}.VfPpkd-WsjYwc{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-sizing:border-box;box-sizing:border-box}.VfPpkd-WsjYwc::after{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-WsjYwc::after{border-color:CanvasText}}.VfPpkd-WsjYwc-OWXEXe-INsAgc::after{border:none}.VfPpkd-aGsRMb{border-radius:inherit;height:100%}.VfPpkd-gBNGNe{position:relative;-moz-box-sizing:border-box;box-sizing:border-box;background-repeat:no-repeat;background-position:center;background-size:cover}.VfPpkd-gBNGNe::before{display:block;content:""}.VfPpkd-gBNGNe:first-child{border-top-left-radius:inherit;border-top-right-radius:inherit}.VfPpkd-gBNGNe:last-child{border-bottom-left-radius:inherit;border-bottom-right-radius:inherit}.VfPpkd-gBNGNe-OWXEXe-BaYisc::before{margin-top:100%}.VfPpkd-gBNGNe-OWXEXe-W3lGp-Clt0zb::before{margin-top:56.25%}.VfPpkd-gBNGNe-bN97Pc{position:absolute;top:0;right:0;bottom:0;left:0;-moz-box-sizing:border-box;box-sizing:border-box}.VfPpkd-EScbFb-JIbuQc{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-sizing:border-box;box-sizing:border-box;position:relative;outline:none;color:inherit;text-decoration:none;cursor:pointer;overflow:hidden}.VfPpkd-EScbFb-JIbuQc:first-child{border-top-left-radius:inherit;border-top-right-radius:inherit}.VfPpkd-EScbFb-JIbuQc:last-child{border-bottom-left-radius:inherit;border-bottom-right-radius:inherit}.VfPpkd-gqIiZe{display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;-moz-box-align:center;align-items:center;-moz-box-sizing:border-box;box-sizing:border-box;min-height:52px;padding:8px}.VfPpkd-gqIiZe-OWXEXe-Vkfede-rJCtOc{padding:0}.VfPpkd-aPoio-c6xFrd,.VfPpkd-aPoio-fuEl3d{display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;-moz-box-align:center;align-items:center;-moz-box-sizing:border-box;box-sizing:border-box}.VfPpkd-aPoio-fuEl3d{color:rgba(0,0,0,.6);-moz-box-flex:1;flex-grow:1;-moz-box-pack:end;justify-content:flex-end}.VfPpkd-aPoio-c6xFrd+.VfPpkd-aPoio-fuEl3d{margin-left:16px;margin-right:0}[dir=rtl] .VfPpkd-aPoio-c6xFrd+.VfPpkd-aPoio-fuEl3d,.VfPpkd-aPoio-c6xFrd+.VfPpkd-aPoio-fuEl3d[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-aPoio{display:-moz-inline-box;display:inline-flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;-moz-box-align:center;align-items:center;-moz-box-sizing:border-box;box-sizing:border-box;-moz-box-pack:center;justify-content:center;cursor:pointer;-moz-user-select:none;user-select:none}.VfPpkd-aPoio:focus{outline:none}.VfPpkd-aPoio-OWXEXe-LgbsSe{margin-left:0;margin-right:8px;padding:0 8px}[dir=rtl] .VfPpkd-aPoio-OWXEXe-LgbsSe,.VfPpkd-aPoio-OWXEXe-LgbsSe[dir=rtl]{margin-left:8px;margin-right:0}.VfPpkd-aPoio-OWXEXe-LgbsSe:last-child{margin-left:0;margin-right:0}[dir=rtl] .VfPpkd-aPoio-OWXEXe-LgbsSe:last-child,.VfPpkd-aPoio-OWXEXe-LgbsSe:last-child[dir=rtl]{margin-left:0;margin-right:0}.VfPpkd-gqIiZe-OWXEXe-Vkfede-rJCtOc .VfPpkd-aPoio-OWXEXe-LgbsSe{-moz-box-pack:justify;justify-content:space-between;width:100%;height:auto;max-height:none;margin:0;padding:8px 16px;text-align:left}[dir=rtl] .VfPpkd-gqIiZe-OWXEXe-Vkfede-rJCtOc .VfPpkd-aPoio-OWXEXe-LgbsSe,.VfPpkd-gqIiZe-OWXEXe-Vkfede-rJCtOc .VfPpkd-aPoio-OWXEXe-LgbsSe[dir=rtl]{text-align:right}.VfPpkd-aPoio-OWXEXe-Bz112c{margin:-6px 0;padding:12px}.VfPpkd-aPoio-OWXEXe-Bz112c:not(:disabled){color:rgba(0,0,0,.6)}.VfPpkd-EScbFb-JIbuQc{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::before,.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::before{transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-FJ5hab::before{transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-FJ5hab::after{top:0;left:0;transform:scale(0);transform-origin:center center}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-FJ5hab::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-FJ5hab::after{animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-FJ5hab::after{animation:mdc-ripple-fg-opacity-out .15s;transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::before,.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::after{top:-50%;left:-50%;width:200%;height:200%}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d .VfPpkd-FJ5hab::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::before,.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-EScbFb-JIbuQc:hover .VfPpkd-FJ5hab::before,.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-FJ5hab::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-FJ5hab::before,.VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-FJ5hab::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-FJ5hab::after{transition:opacity .15s linear}.VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-FJ5hab::after{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab{-moz-box-sizing:content-box;box-sizing:content-box;height:100%;overflow:hidden;left:0;pointer-events:none;position:absolute;top:0;width:100%}.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::after,.VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):focus::after{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:5px double transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::after,.VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):focus::after{border-color:CanvasText}}.KC1dQ{border-radius:8px;background-color:#fff;border-width:0;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15)}.KC1dQ .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Usd1Ac{border-radius:8px;background-color:#fff;border:1px solid rgb(218,220,224);box-shadow:none}.Usd1Ac .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Si6A0c{position:absolute;left:0;top:0;width:100%;height:100%;outline:none}.MONpF{background:rgb(206,234,214);border-radius:52px;color:rgb(13,101,45);line-height:20px;margin-left:1rem;padding:0 .375rem;text-align:center;font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.bg6sud{margin-bottom:-0.5rem}.xtiq3{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:wrap;flex-wrap:wrap}.N33kHb{margin-left:1.5rem;padding-top:1rem}.UJYYgf{margin-right:0.5rem}.Lqr2e{background-position:center center;background-repeat:no-repeat;background-size:contain;flex-shrink:1;height:23.75rem;margin-bottom:1.875rem;max-height:15rem;width:90%}.KUqHO{box-sizing:border-box;justify-content:flex-start;padding-top:7.5rem;text-align:center}.KUqHO h1,.KUqHO h2{margin-bottom:1.5rem}.ZLgLX{align-items:center;box-sizing:border-box;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:2rem 1rem 1.5rem;text-align:center;width:18.75rem}.ZLgLX .Lqr2e{height:7.375rem}@media (max-height:35.5em){.UrFp8e .Lqr2e{height:40%;margin-bottom:0.5rem}}.WagS8{margin-bottom:0}.hcjKL{position:absolute;right:0.3125rem;top:0.3125rem}.GqugBc{height:4.375rem;position:relative;left:1.9375rem}.nt2KVb{width:11.25rem}.nfX1Z{margin:0.5rem 0.5rem 0}.CJZRbc{margin-top:-1rem}.Vo9Zre{display:inline-block}.Vo9Zre h1{margin-left:1.5rem;margin-top:3.375rem}.Vo9Zre .EIsTbe{display:inline-block;margin-left:1.5rem;margin-top:1.5rem}.Vo9Zre .nQIsGb{margin:0 auto;max-width:15rem}.CxlSNe{color:rgb(95,99,104)}.CxlSNe:not(:empty){padding-left:16px}.nHTcze{display:-moz-box;display:flex;-moz-box-align:center;align-items:center}.R7HDBc{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400}@media not (min-width:600px){.R7HDBc{display:none}}@media (min-width:600px){.nHTcze{display:none}}.cBtBT{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-flex:1;flex-grow:1;min-width:0}.R2KREf{-moz-box-align:center;align-items:center;background:#fff;display:-moz-box;display:flex;height:48px;-moz-box-pack:justify;justify-content:space-between;min-width:0;padding-left:16px}.TlWbF,.EgTw4e .qRUolc{border-bottom:1px solid rgba(0,0,0,.12)}.UE04Dc{height:24px;padding-right:16px;width:24px}.qSxFt{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-flex:1;flex-grow:1;min-width:0}.pEh7df{margin-left:8px}.dj7Enb .X1clqd .R2KREf{margin:-16px}.dj7Enb .qRUolc .R2KREf{margin:-18px -24px -16px}.dj7Enb .qRUolc .pPQgvf{margin:0}.dj7Enb .wnIM7{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;padding:0}.EgTw4e{height:80%}.T9Iutc{margin-right:8px}@media (max-width:600px){.EgTw4e{max-width:none;width:100%}}@media not all and (max-width:600px){.EgTw4e{max-width:1600px;width:90%}}.gqPc8{border-width:0;-moz-box-sizing:border-box;box-sizing:border-box;-moz-box-flex:1;flex-grow:1}.tthERc{position:absolute;border:none;width:100%;height:calc(100vh - 4.0625rem)}.X65jac{margin-bottom:1rem}.zxFw5d{margin-bottom:1.5rem}.Elz9Mb{-moz-box-flex:1 1 100%;flex:1 1 100%;overflow:hidden}.BuI5lb{margin-right:1rem}.PtHAPb{margin-right:0.375rem}.E5l1S{-moz-box-flex:none;flex:none}.E5f6Vd{border-top:0.0625rem solid #e0e0e0;margin:0 -1.5rem 1.5rem}.f2YrEb{padding-bottom:0.5rem}.ipmZkd{margin-bottom:.5rem}.FLgDTb{padding:1.5rem;margin-bottom:2rem}.NXcbkc{margin-top:1rem}.NGiYh.NGiYh.NGiYh.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-pafCAf{fill:transparent}.NGiYh.NGiYh.NGiYh.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-pafCAf{fill:transparent}.NGiYh.NGiYh.NGiYh.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled .VfPpkd-pafCAf{fill:transparent}.NGiYh.NGiYh.NGiYh.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-pafCAf{fill:transparent}.io4oZb{margin-bottom:1rem}.UiyBvb .io4oZb .JYB4b{margin-bottom:1rem;padding:0}.qXTVSe{margin:0.5rem 0}.uQNHvf.uQNHvf{height:32px;margin-right:0.5rem;width:32px}.EfLcNb{margin-bottom:1rem}.gJJVDc{height:3rem;width:3rem}.jkutNd{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.ESVbeb,.W9d6ec{color:rgb(95,99,104);margin:.5rem}.ESVbeb{width:15rem}.j2VD8e{text-align:center}.QIo6w{margin-top:.75rem;text-align:right;width:15rem}.a2Umne{margin-top:.5rem}.ljCLXb{-moz-box-align:center;align-items:center;background:white;bottom:0;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;left:0;padding-top:1rem;position:fixed;right:0;top:4rem}.Pp6l6e{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;margin:1rem}.FomsT{display:block;margin:.75rem;width:15rem}.kwpuYb{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.FomsT .oJeWuf{-moz-box-align:center;align-items:center}.FomsT .Qks78e{height:2.5rem}.FomsT .JtDYBc{margin-right:.5rem}.kX9r6c{margin:.5rem auto;max-width:25rem;padding:.5rem}.TLI4vb{margin-right:1rem}.KUHggb{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.n5lRPb{margin-top:.25rem}.a3O8K{margin:1.5rem 0}.m9odT{margin-top:.75rem;text-align:right}.LDr2ne{border-bottom:0.0625rem solid #e0e0e0;border-top:0.0625rem solid #e0e0e0;margin:0 -1.5rem 1rem -1.5rem;padding:1rem 1.5rem}.xS7jB{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:space-between}.D9l13b{color:rgba(0,0,0,.549);margin:0.5rem 0 0.25rem 0}.rLpHLd{max-width:none}.cdsSCb{display:inline-block;border-bottom:1px solid currentColor;line-height:1em;vertical-align:top;width:1.5em}.regK8{-moz-box-align:stretch;align-items:stretch;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.UHsoGd.UHsoGd{width:auto}.UHsoGd .zHQkBf{padding:8px 0 8px 8px;text-align:right;color:inherit;font-family:inherit;font-size:inherit;font-weight:inherit;letter-spacing:inherit;line-height:inherit}.UHsoGd .MQL3Ob{flex-shrink:0;max-width:40%;padding-left:0;padding-right:8px}.hbAdzc{white-space:nowrap}.fJiTAb .RxsGPe{font-size:.1rem;height:.1rem;line-height:1;opacity:.001;overflow:hidden;position:absolute;width:.1rem}.HgKLRe .zHQkBf{color:inherit;font-family:inherit;font-size:inherit;font-weight:inherit;letter-spacing:inherit;line-height:inherit}.HgKLRe:not(.fvAYpc) .zHQkBf{text-align:right}.HgKLRe.fvAYpc .zHQkBf{text-align:right}.YeoM1d{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;height:100%;white-space:nowrap}.HgKLRe .MQL3Ob{flex-shrink:0;max-width:40%}.HgKLRe:not(.fvAYpc) .MQL3Ob{padding-left:0}.HgKLRe.fvAYpc .MQL3Ob{direction:ltr;padding-left:0}.DAadud .zHQkBf{padding:8px}.DAadud:not(.fvAYpc) .zHQkBf{padding-right:0}.DAadud.fvAYpc .zHQkBf{padding-right:0}.DAadud:not(.fvAYpc) .MQL3Ob{padding-right:8px}.DAadud.fvAYpc .MQL3Ob{padding-right:8px}.E9XmEd{-moz-box-align:stretch;align-items:stretch;display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.E9XmEd .jlfrG{-moz-box-flex:0;-moz-box-flex:0 0 200px;flex:0 0 200px;min-height:150px;width:200px}.E9XmEd .jlfrG:not(:last-child){margin-right:8px}.Q35ysf{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.Q35ysf .jlfrG{flex-shrink:0}.Q35ysf .jlfrG:not(:last-child){margin-bottom:8px}.jlfrG{color:#3c4043;display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;overflow-y:hidden;position:relative}.lnAGpc{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1;-moz-box-flex:1 1 auto;flex:1 1 auto;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;outline:none;overflow-x:hidden;overflow-y:auto;padding:8px 16px;position:relative}.jlfrG:before,.jlfrG:after{content:"";height:8px;left:0;position:absolute;right:0}.jlfrG:before{background:linear-gradient(to bottom,#fff,transparent);top:0;z-index:1}.jlfrG:after{background:linear-gradient(to top,#fff,transparent);bottom:0}.E9XmEd .jlfrG{max-height:216px}.Q35ysf .jlfrG{max-height:166px}.VBYA0c{-moz-box-align:start;align-items:flex-start;display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-shrink:0;margin-bottom:8px}.ILZUr{-moz-box-flex:1;box-flex:1;flex-grow:1;margin-right:8px}.iaDxJf{font-style:italic;text-align:end}.pN6IZc{flex-shrink:0}.rhVLBd{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.OK1tJe:not(:last-child){margin-right:4px}.OK1tJe{background-color:#f1f3f4;-moz-border-radius:2px;border-radius:2px;-moz-box-flex:1;-moz-box-flex:1 1 auto;flex:1 1 auto;height:24px;outline:none}.R5iLrf.KKjvXb .lnAGpc,.R5iLrf.KKjvXb.OK1tJe{outline:1px dashed transparent}.R5iLrf.u3bW4e .lnAGpc,.R5iLrf.u3bW4e.OK1tJe{outline:1px solid transparent}.R5iLrf.yXgmRe:hover{cursor:pointer}.R5iLrf.u3bW4e,.R5iLrf.yXgmRe:hover{background-color:#e8eaed}.jlfrG.u3bW4e:before,.jlfrG.yXgmRe:hover:before{background:linear-gradient(to bottom,#e8eaed,transparent)}.jlfrG.u3bW4e:after,.jlfrG.yXgmRe:hover:after{background:linear-gradient(to top,#e8eaed,transparent)}.R5iLrf.KKjvXb{background-color:#1a73e8;color:#fff}.jlfrG.KKjvXb:before{background:linear-gradient(to bottom,#1a73e8,transparent)}.jlfrG.KKjvXb:after{background:linear-gradient(to top,#1a73e8,transparent)}.R5iLrf.KKjvXb.u3bW4e,.R5iLrf.KKjvXb.yXgmRe:hover{background-color:#1967d2}.jlfrG.KKjvXb.u3bW4e:before,.jlfrG.KKjvXb.yXgmRe:hover:before{background:linear-gradient(to bottom,#1967d2,transparent)}.jlfrG.KKjvXb.u3bW4e:after,.jlfrG.KKjvXb.yXgmRe:hover:after{background:linear-gradient(to top,#1967d2,transparent)}.NBQ1Tb.noVAQc .UGEHab,.NBQ1Tb:not(.noVAQc) .cU5Ufe{display:none}.v2RmYb{display:-moz-box;display:flex}.i8ebQe{-moz-box-align:stretch;align-items:stretch;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.stS1kf{padding:4px 4px 4px 16px}.FMomcc .Fxmcue{text-align:start}.mcDcFb,.FMomcc .snByac{overflow:hidden}.jcygrd{flex-shrink:0;margin-right:4px}.jjKzBb{margin-right:8px}.hlKmZb{width:80px}.o1Okpe{margin-left:4px}.gXJ4Pb{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.UjXaMc{padding:0 16px 16px 16px}.ZtfTEf{margin:4px 24px 8px;text-align:end}.rjqfkb{display:-moz-box;display:flex;overflow-x:auto;overflow-y:hidden}.yxqL6,.tMKXJb{-moz-box-sizing:border-box;box-sizing:border-box;padding:0 16px 16px 16px}.yxqL6{width:300px}.bHR9hf{-moz-box-align:stretch;align-items:stretch;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.aVdG0e{margin-right:5px;margin-bottom:8px}.oPshk{margin-left:11px}.oPshk.Lm9w4d .gWQ8we,.oPshk:not(.Lm9w4d) .ZJxgub{display:none}.E7ZeX{-moz-box-align:stretch;align-items:stretch;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.OK63Pb:not(:last-child){border-bottom:1px solid rgba(0,0,0,.12)}.Z3wmOd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.AgnJoc{font-weight:400}.nl5VRd{margin-bottom:1rem;position:relative}@media (max-width:30em){.nl5VRd{margin-bottom:0.5rem}}.N5dSp{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-bottom:0.25rem}.I0naMd{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:1.75rem;margin-left:0.5rem}.W4hhKd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:space-between;padding-bottom:0.5rem}@media (max-width:30em){.W4hhKd{flex-direction:column}}.CzuI5c:not(:empty){-moz-flex-wrap:wrap;flex-wrap:wrap;margin-bottom:0.5rem;margin-right:1rem;overflow:hidden}.fOvfyc{overflow:hidden;word-wrap:break-word}.rec5Nb{-moz-flex-wrap:wrap;flex-wrap:wrap;margin-bottom:0.5rem}.DwLQSc{margin:0 0.25rem}.DwLQSc:first-of-type,.DwLQSc:last-of-type{display:none}.Wa3mee{margin-bottom:0.5rem}.nGi02b{margin-bottom:1rem;overflow:hidden;word-wrap:break-word}.tWdbMc{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:wrap;flex-wrap:wrap;justify-content:space-between;padding:0.5rem 1rem}.pzyQle{-moz-box-flex:1 0 auto;flex:1 0 auto;justify-content:flex-end}.P47N4e{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;margin-right:1rem}.P47N4e.P47N4e{height:2.375rem;width:2.375rem}.fJ1Vac{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;padding:1.25rem 1.5rem 1.5rem 1.5rem}@media (max-width:30em){.fJ1Vac{padding:0.25rem 0.5rem 0.5rem 0.5rem}}.EE538{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-flex:1 1 auto;flex:1 1 auto;flex-direction:column;max-width:47.5rem;min-width:0}.BiaLW{-moz-box-flex:0 0 auto;flex:0 0 auto;margin-left:2rem;max-width:18.75rem;width:18.75rem}.kwWsO{padding-bottom:0.5rem}.ar1wE .eqqrO,.ySjuvd .eqqrO{border-top:0.125rem solid #e8eaed}.lq45g{padding-top:1rem}.AJFihd{padding:1.5rem}.Dy8Cxc{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:wrap;flex-wrap:wrap;justify-content:space-between;margin-bottom:0.5rem}.KI1A1e{text-align:right}.P2wHlc{border-bottom:0.0625rem solid #e0e0e0;margin-bottom:1rem}.B2pRjc{margin:2rem 0;text-align:center}.IPGLSb{align-items:stretch;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.cYYbdd{margin-bottom:1rem}.XgQDH{padding-bottom:0.5rem;padding-top:0.5rem}.QxGMXc{margin:1rem 1.5rem 0 1.5rem}.uGeUQe{margin-left:-0.5rem}.Epqnjf{margin:0 1.25rem}.lLBkgb:not(:empty){margin-bottom:1rem}.hjqfGd{padding-bottom:1rem}@media (max-width:30em){.hjqfGd{padding-bottom:0}}.sGidkc .kCI6s{width:8rem}.uyN3Kb .kCI6s{width:10rem}.sGidkc .RSOxzc,.uyN3Kb .RSOxzc{width:100%}.CNB7te{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:100%;justify-content:space-between;line-height:1}.FEOARd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.f5Kwpe{box-sizing:border-box;flex-shrink:0;padding-left:4.25rem;padding-right:1.5rem;width:28rem}.wvJNcc{box-sizing:border-box;flex-shrink:0;padding:0.75rem 1rem 0.75rem 1.5rem;width:28rem}.UumJte{margin-right:1rem;flex-shrink:0}.bCoXYd{width:1.5rem}.CNB7te>:last-child{flex-shrink:0;margin-right:1rem}.wvJNcc>:last-child{flex-shrink:0;margin-left:auto}@media (max-width:61.25em){.f5Kwpe,.wvJNcc{box-flex:1;flex-grow:1;flex-shrink:1;width:auto;padding-right:0}.wvJNcc>:last-child{margin-right:1rem}.CNB7te>:last-child{margin-right:1.5rem}}@media (max-width:30em){.f5Kwpe>.Nmpzvc{-moz-box-flex:1 11 0.5rem;flex:1 11 0.5rem}.CNB7te>:last-child{margin-right:1rem}}@media (max-width:25em){.f5Kwpe{padding-left:1rem}.UumJte{margin-right:0.5rem}.CNB7te>:last-child{margin-right:0}}.hLVkAc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;max-width:100%}.j6EwUd{background:#e8eaed;-moz-border-radius:0.25rem;border-radius:0.25rem;gap:0.5rem;overflow:hidden;padding:0.25rem 0.5rem}.jPglrc{height:1.5rem;width:1.5rem}.B71iyf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;min-width:0}.Q7YAVc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.dWdaJc{text-overflow:ellipsis;overflow:hidden;white-space:nowrap}.Jc6qh{border-color:rgb(60,64,67)}.oqnjOc table{border-collapse:collapse;position:relative;width:100%}.fWM9Tb{height:3rem}.TAjiIf a{align-items:center;color:inherit;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:100%;text-decoration:none}.TJtJXb .TAjiIf a:focus .ZcoGnf,.TJtJXb .TAjiIf a:hover .ZcoGnf,.tYQn5c .TAjiIf a:focus,.tYQn5c .TAjiIf a:hover,.DC55n .TAjiIf a:focus .MNAqQb,.DC55n .TAjiIf a:hover .MNAqQb{text-decoration:underline}.oqnjOc td{height:4rem;padding:0;padding-left:1.5rem}.oqnjOc td.TAjiIf{max-width:0;overflow:hidden;padding-right:1rem}.oqnjOc td.TAjiIf:last-child{padding-right:1.5rem}.JlndIc{overflow:hidden}.pNoxUe{width:1.25rem}.LiCTz{width:100%}.Fk0vXe{width:8.25rem}.TJtJXb .TAjiIf .vUBwW{margin-right:1rem}.uGg1kd,.wpvRpe{position:relative}.oWYiGe{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-flow:column wrap;gap:0.5rem;margin:0.5rem 0.5rem 0.5rem 0}.VUdUqf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-flow:column wrap;gap:0.5rem;margin:0.75rem 0.5rem 0.75rem 0}.hn7AEc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:wrap;flex-wrap:wrap;justify-content:space-between;gap:0.5rem}.RAboLe{margin-right:0}.nTrDbc .uGg1kd{padding-left:4.25rem}.nTrDbc .wpvRpe{padding-left:2.5rem}.DC55n td{background:white;border-top:0.0625rem solid #e0e0e0;border-bottom:0.0625rem solid #e0e0e0}.DC55n .tkmmwb{margin-right:1rem}.oqnjOc td.Fk0vXe{border-left:0.0625rem solid #e0e0e0;padding:0}.TJtJXb:hover td,.tYQn5c:hover td,.DC55n:hover td{background:#f5f5f5}.aSjeL.aSjeL td{background:#f5f5f5}.gyaw1d .oqnjOc .oFj0xc{cursor:pointer}.CgLVWe.CgLVWe{height:100%;overflow:hidden}.CgLVWe .T4LgNb,.CgLVWe .kFwPee:not(.OOnEBd),.DReKqd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;height:100%;overflow:hidden}.BQ5ILd{border-bottom:0.0625rem solid #e0e0e0;flex-shrink:0;height:4rem}.mthue{align-items:stretch;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;box-flex:1;flex-grow:1;overflow:hidden}.lBRpOc{flex-shrink:0;overflow:auto;position:relative;width:28rem}.a4YS1c{border-left:0.0625rem solid #e0e0e0;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:1;flex-grow:1;overflow:hidden}@media (max-width:61.25em){.lBRpOc{box-flex:1;flex-grow:1;flex-shrink:1;overflow-x:hidden;overflow-y:visible;width:auto}.a4YS1c{border-left:none}}@media not all and (max-width:61.25em){.jBWfpf.jBWfpf{display:none}}@media (max-width:61.25em){.Alnfpc.Alnfpc{display:none}}.CcC9kf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;box-flex:1;flex-grow:1;overflow:auto}.CcC9kf>*{flex-shrink:0}.ALvsPd{padding:1.5rem;padding-bottom:0}.xPSjRb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:space-between;margin-bottom:1rem}.kHjrfc:not(:empty){margin-top:1rem}@media not all and (max-width:30em){.DReKqd .yHjGtf:nth-child(1),.DReKqd .yHjGtf:nth-child(2){border-left:none;padding-left:0}}.OFjtS{height:3rem}.XsISn{margin:0.5rem 0 1.5rem 1rem}.g5FCDc{border-top:0.0625rem solid #e0e0e0;overflow:hidden}@media (max-width:61.25em){.gyaw1d .BQ5ILd,.gyaw1d .lBRpOc{display:none}}.I2pI{font-size:0.875rem;margin-right:1rem}.iq6Osb{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding-bottom:4rem;padding-top:4rem}@media (max-width:40em){.iq6Osb{padding-top:1.5rem}}@media not all and (max-width:40em){.YXGmid{margin-top:4.375rem}}.YXGmid .BgnnGb{height:9.375rem}.yfjJPb{margin-bottom:0.5rem;margin-top:1.5rem}.jFNEDb{text-align:center;max-width:17.5rem}.MHxtic{margin:0 1.5rem;padding:1rem 0}.MHxtic:not(:last-child){border-bottom:0.0625rem solid #e0e0e0}@media (max-width:48.75em){.MHxtic{margin:0 1.5rem}.MHxtic:first-child{margin-top:-1rem}.MHxtic:last-child{margin-bottom:-1rem}}@media (max-width:30em){.MHxtic{margin:0 1rem}}@media not all and (max-width:30em){.MHxtic:hover{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);border-radius:0.5rem;margin-left:0;margin-right:0;overflow:hidden;padding-left:1.5rem;padding-right:1.5rem}}.MHxtic:focus-within{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);border-radius:0.5rem;margin-left:0;margin-right:0;overflow:hidden;padding-left:1.5rem;padding-right:1.5rem}@media (max-width:30em){.MHxtic:focus-within{padding-left:1rem;padding-right:1rem}}.nUg0Te{text-decoration:none;box-flex:1;flex-grow:1;min-width:0}.mh4Cme{align-self:start;-moz-border-radius:50%;border-radius:50%;flex-shrink:0;height:2.25rem;width:2.25rem}.ZHEgO{opacity:0.26}.il4hc,.XQMoHb{-moz-box-flex:1;flex:1;min-width:0}.il4hc{padding-left:1rem}.XQMoHb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}@media (max-width:30em){.XQMoHb{flex-direction:column}.e5iAof{padding-left:3.25rem;padding-top:1rem}}@media not all and (max-width:30em){.XQMoHb{flex-direction:row}}.tGZ0W{align-self:center;margin-left:1.5rem;text-align:right}@media (max-width:40em){.tGZ0W{align-self:start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}}.iiWxqc{margin-top:0.75rem}.mN0Vkf{color:#9aa0a6}.SBb9Ed{font-style:italic;text-align:right}.y9bEQb{-moz-box-flex:1;flex:1;min-width:0}.y9bEQb>*:not(:last-child){margin-bottom:0.25rem}.LKqFXc{border-top:0.0625rem solid #e0e0e0;margin:0 1.5rem;padding-top:1rem}@media (max-width:48.75em){.LKqFXc{margin-top:1rem}}.x39Mke{padding-left:1.5rem;padding-bottom:1.5rem}@media (max-width:48.75em){.x39Mke{padding-left:0}}@media (max-width:30em){.x39Mke{padding:1rem 0.5rem}}.fzV7Xc{margin-bottom:1.5rem}.NLc53c{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.125rem;font-weight:400;letter-spacing:0;line-height:1.5rem;color:#3c4043;padding-left:1.5rem;margin-bottom:1rem}.YH8M6e{margin-bottom:0.25rem}.mQtmBc{padding-right:1.5rem}.B0fUvb{color:#9aa0a6}@media not all and (max-width:48.75em){.XAGGOd{margin-right:-0.5rem}}@media (max-width:30em){.NLc53c{padding-left:1rem}.NLc53c:first-child{margin-top:1rem}.hmNEpf{align-self:start;padding-top:0.25rem}}.e0Cfsd{border-radius:1.5rem;-moz-box-sizing:border-box;box-sizing:border-box;height:35rem;max-width:43.75rem;position:relative;width:100%}.RMDLeb{height:100%}.eNJEwd,.i5sehe,.kox42c{-moz-box-sizing:border-box;box-sizing:border-box;height:100%;overflow:hidden;width:100%}.i5sehe.i5sehe,.l73pue .Jj5MRb.kox42c{overflow-y:auto}.i5sehe,.kox42c{-moz-box-align:center;align-items:center;background-color:#fff;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;left:0;padding:2rem;position:absolute;top:0}.i5sehe{opacity:1;z-index:1}@media (max-width:40rem){.e0Cfsd{border-radius:0;bottom:0;box-shadow:none;height:100%;left:0;max-width:100%;overflow:auto;position:fixed;right:0;top:0;width:100%}}@media (max-width:30rem){.eNJEwd{padding:.5rem}.NZ9wdc{padding:1rem 1rem 0 1rem}}.NZ9wdc{align-self:stretch;-moz-box-align:center;align-items:center;background-color:rgb(248,249,250);-moz-box-sizing:border-box;box-sizing:border-box;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;height:19.625rem;margin:-2rem -2rem 0 -2rem;padding:2rem 2rem 0 2rem}.i5sehe.TfD4bb{margin-left:-100%;opacity:0;transition:margin-left .5s cubic-bezier(.4,0,.2,1),opacity .5s cubic-bezier(.4,0,.2,1)}.i5sehe.TfD4bb .O0WRkf{visibility:hidden}.bQEkKf,.clp6rf{text-align:center;max-width:26.5625rem}.SVDBnd{margin-top:1.5rem}.i5sehe .aP3ZPb{bottom:0;position:absolute}.rsGJMc{max-width:100%}.GHskLb{padding:0 .5rem;position:relative}.LeM6cb{margin-top:-1rem;margin-bottom:2rem;text-align:center;width:100%}.A0jDm{background-color:white;display:block;height:18rem}.A0jDm{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15)}.A0jDm.A0jDm:not(.RDPZE){border:none}.lLzY8b:not(:first-child){margin-left:1.5rem}@media (max-width:30rem){.lLzY8b:not(:first-child){margin-left:.5rem}}.A0jDm.RDPZE .snByac>*:not(.aP3ZPb){opacity:.37}.A0jDm.A0jDm .Fxmcue{display:block;height:100%;padding:0}.A0jDm .snByac{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;line-height:1.75rem;-moz-box-align:center;align-items:center;color:rgb(60,64,67);display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;padding:2rem}.zBlW2d{max-width:100%;width:10.5rem;margin-bottom:1.5rem}.A0jDm .aP3ZPb{left:0;position:absolute;right:0;top:0;z-index:1}.EDId0c{position:relative}.nhh4Ic{position:absolute;left:0;right:0;top:0;z-index:1;pointer-events:none}.nhh4Ic[data-state=snapping],.nhh4Ic[data-state=cancelled]{-moz-transition:transform 200ms;transition:transform 200ms}.MGUFnf{display:block;width:28px;height:28px;padding:15px;margin:0 auto;transform:scale(0.7);background-color:#fafafa;border:1px solid #e0e0e0;-moz-border-radius:50%;border-radius:50%;-moz-box-shadow:0 2px 2px 0 rgba(0,0,0,.2);box-shadow:0 2px 2px 0 rgba(0,0,0,.2);-moz-transition:opacity 400ms;transition:opacity 400ms}.nhh4Ic[data-state=resting] .MGUFnf,.nhh4Ic[data-state=cooldown] .MGUFnf{transform:scale(0);-moz-transition:transform 150ms;transition:transform 150ms}.nhh4Ic .LLCa0e{stroke-width:3.6px;-moz-transform:translateZ(1px);transform:translateZ(1px)}.nhh4Ic[data-past-threshold=false] .LLCa0e{opacity:.3}.rOhAxb{fill:#4285f4;stroke:#4285f4}.A6UUqe{display:none;stroke-width:3px;width:28px;height:28px}.tbcVO{width:28px;height:28px}.bQ7oke{position:absolute;width:0;height:0;overflow:hidden}.A6UUqe.qs41qe{animation-name:quantumWizSpinnerRotate;animation-duration:1568.63ms;animation-iteration-count:infinite;animation-timing-function:linear;display:inline-block}.A6UUqe.SdoWjb{display:inline-block}.A6UUqe.qs41qe .ceIWpc{stroke:none;fill:none}.A6UUqe.sf4e6b .qjUCkf{stroke-width:0}.qjUCkf{-moz-transition:stroke-width 400ms;transition:stroke-width 400ms;transform-origin:14px 14px;stroke-dasharray:58.9 58.9;stroke-dashoffset:58.9;fill:none;-moz-transform:rotate(0deg);transform:rotate(0deg)}.A6UUqe.SdoWjb .qjUCkf{transition-duration:0}.A6UUqe.iPwZeb .qjUCkf{animation-delay:-466ms,-466ms,-466ms}.A6UUqe.qs41qe .qjUCkf{animation-name:quantumWizSpinnerFillUnfill,quantumWizSpinnerRot,quantumWizSpinnerColors;animation-duration:1333ms,5332ms,5332ms;animation-iteration-count:infinite,infinite,infinite;animation-timing-function:cubic-bezier(0.4,0,0.2,1),steps(4),linear;animation-fill-mode:forwards}@keyframes quantumWizSpinnerRotate{0%{-moz-transform:rotate(0deg);transform:rotate(0deg)}to{-moz-transform:rotate(360deg);transform:rotate(360deg)}}@keyframes quantumWizSpinnerFillUnfill{0%{stroke-dashoffset:58.8}50%{stroke-dashoffset:0}to{stroke-dashoffset:-58.4}}@keyframes quantumWizSpinnerRot{0%{-moz-transform:rotate(0deg);transform:rotate(0deg)}to{-moz-transform:rotate(-360deg);transform:rotate(-360deg)}}@keyframes quantumWizSpinnerColors{0%{stroke:#4285f4}18%{stroke:#4285f4}25%{stroke:#db4437}43%{stroke:#db4437}50%{stroke:#f4b400}68%{stroke:#f4b400}75%{stroke:#0f9d58}93%{stroke:#0f9d58}to{stroke:#4285f4}}.zpf6Qc{height:100%;overflow-y:auto}.zpf6Qc .fkiogf{display:block}.zpf6Qc .dNuvt{-moz-box-align:center;align-items:center;-moz-box-sizing:border-box;box-sizing:border-box;display:-moz-box;display:flex;-moz-box-pack:center;justify-content:center;padding:8px;width:100%}.thP79c{-moz-user-select:none;-moz-transition:background-color .1s ease;transition:background-color .1s ease;align-items:center;box-sizing:border-box;cursor:pointer;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;font-weight:500;min-height:48px;line-height:20px;outline:none;overflow:hidden;padding:12px 16px;position:relative}.thP79c.fEAHmc{padding:8px 16px}.thP79c.C2k2wf{align-items:flex-start}.sU5zjc,.Yrzgvb{-moz-border-radius:50%;border-radius:50%;height:40px;width:40px}.p8ihof{margin-right:16px}.OeTIXd{min-width:0}.thP79c:hover{background-color:rgba(32,33,36,0.039)}.lRaOFf[aria-selected="true"]{background-color:rgba(32,33,36,0.078)}.lRaOFf[aria-selected="true"]:hover{background-color:rgba(32,33,36,0.102)}.thP79c:focus,.lRaOFf[aria-selected="true"]:focus{background-color:rgba(32,33,36,0.122)}.thP79c:focus:hover{background-color:rgba(32,33,36,0.157)}.thP79c.qs41qe,.thP79c.qs41qe:focus,.thP79c.qs41qe:hover{background-color:rgba(32,33,36,0.157)}.thP79c.RDPZE,.thP79c.RDPZE:hover,.thP79c.RDPZE:focus{background-color:transparent;color:rgba(0,0,0,.26)}.nNi7jd.C2k2wf,.n0MHff.C2k2wf{padding:16px}.DRS7P,.eL4rW{overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.p9A2Ge{overflow:hidden;text-overflow:ellipsis;white-space:nowrap;color:rgba(0,0,0,.54);font-size:14px;line-height:20px}.thP79c.RDPZE .p9A2Ge{color:rgba(0,0,0,.12)}.Sg7FOe{-moz-transform:translate(-50%,-50%) scale(0);transform:translate(-50%,-50%) scale(0);-moz-transition:opacity .3s ease;transition:opacity .3s ease;background-size:cover;left:0;opacity:0;pointer-events:none;position:absolute;top:0}.thP79c.qs41qe .Sg7FOe{transition:-webkit-transform 0.3s cubic-bezier(0,0,0.2,1);transition:transform 0.3s cubic-bezier(0,0,0.2,1);-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2);opacity:1}.thP79c.j7nIZb .Sg7FOe{-moz-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2)}.thP79c .Sg7FOe{background-image:radial-gradient(circle farthest-side,rgba(32,33,36,0.078),rgba(32,33,36,0.078) 80%,rgba(32,33,36,0) 100%)}.eL4rW{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.KL4X6e{background:#eee;bottom:0;left:0;opacity:0;position:absolute;right:0;top:0}.TuA45b{opacity:.8}.VfPpkd-YAxtVc{background-color:#333333}.VfPpkd-gIZMF{color:rgba(255,255,255,.87)}.VfPpkd-YAxtVc{min-width:344px}@media (max-width:344px),(max-width:480px){.VfPpkd-YAxtVc{min-width:100%}}.VfPpkd-YAxtVc{max-width:672px}.VfPpkd-YAxtVc{box-shadow:0 3px 5px -1px rgba(0,0,0,.2),0 6px 10px 0 rgba(0,0,0,.14),0 1px 18px 0 rgba(0,0,0,.12)}.VfPpkd-YAxtVc{border-radius:4px;border-radius:var(--mdc-shape-small,4px)}.VfPpkd-Ng57nc{display:none;position:fixed;right:0;bottom:0;left:0;-moz-box-align:center;align-items:center;-moz-box-pack:center;justify-content:center;-moz-box-sizing:border-box;box-sizing:border-box;pointer-events:none;-webkit-tap-highlight-color:rgba(0,0,0,0)}.VfPpkd-Ng57nc-OWXEXe-uGFO6d,.VfPpkd-Ng57nc-OWXEXe-FNFY6c,.VfPpkd-Ng57nc-OWXEXe-FnSee{display:-moz-box;display:flex}.VfPpkd-Ng57nc-OWXEXe-FNFY6c .VfPpkd-gIZMF,.VfPpkd-Ng57nc-OWXEXe-FNFY6c .VfPpkd-M6tBBc{visibility:visible}.VfPpkd-YAxtVc{padding-left:0;padding-right:8px;display:-moz-box;display:flex;-moz-box-align:center;align-items:center;-moz-box-pack:start;justify-content:flex-start;-moz-box-sizing:border-box;box-sizing:border-box;transform:scale(.8);opacity:0}.VfPpkd-YAxtVc::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-YAxtVc::before{border-color:CanvasText}}[dir=rtl] .VfPpkd-YAxtVc,.VfPpkd-YAxtVc[dir=rtl]{padding-left:8px;padding-right:0}.VfPpkd-Ng57nc-OWXEXe-FNFY6c .VfPpkd-YAxtVc{transform:scale(1);opacity:1;pointer-events:auto;transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),transform .15s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-Ng57nc-OWXEXe-FnSee .VfPpkd-YAxtVc{transform:scale(1);transition:opacity 75ms 0ms cubic-bezier(.4,0,1,1)}.VfPpkd-gIZMF{padding-left:16px;padding-right:8px;width:100%;-moz-box-flex:1;flex-grow:1;-moz-box-sizing:border-box;box-sizing:border-box;margin:0;visibility:hidden;padding-top:14px;padding-bottom:14px}[dir=rtl] .VfPpkd-gIZMF,.VfPpkd-gIZMF[dir=rtl]{padding-left:8px;padding-right:16px}.VfPpkd-gIZMF::before{display:inline;content:attr(data-mdc-snackbar-label-text)}.VfPpkd-M6tBBc{display:-moz-box;display:flex;flex-shrink:0;-moz-box-align:center;align-items:center;-moz-box-sizing:border-box;box-sizing:border-box;visibility:hidden}.VfPpkd-IkaYrd+.VfPpkd-TolmDb{margin-left:8px;margin-right:0}[dir=rtl] .VfPpkd-IkaYrd+.VfPpkd-TolmDb,.VfPpkd-IkaYrd+.VfPpkd-TolmDb[dir=rtl]{margin-left:0;margin-right:8px}.VfPpkd-Ng57nc{z-index:8;margin:8px}.VfPpkd-Ng57nc-OWXEXe-eu7FSc .VfPpkd-gIZMF{padding-left:16px;padding-right:8px;padding-bottom:12px}[dir=rtl] .VfPpkd-Ng57nc-OWXEXe-eu7FSc .VfPpkd-gIZMF,.VfPpkd-Ng57nc-OWXEXe-eu7FSc .VfPpkd-gIZMF[dir=rtl]{padding-left:8px;padding-right:16px}.VfPpkd-Ng57nc-OWXEXe-eu7FSc .VfPpkd-YAxtVc{-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-align:start;align-items:flex-start}.VfPpkd-Ng57nc-OWXEXe-eu7FSc .VfPpkd-M6tBBc{align-self:flex-end;margin-bottom:8px}.VfPpkd-Ng57nc-OWXEXe-M1Soyc{-moz-box-pack:start;justify-content:flex-start}.VfPpkd-gIZMF{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit)}.VfPpkd-IkaYrd:not(:disabled){color:#bb86fc}.VfPpkd-IkaYrd .VfPpkd-Jh9lGc::before,.VfPpkd-IkaYrd .VfPpkd-Jh9lGc::after{background-color:#bb86fc;background-color:var(--mdc-ripple-color,#bb86fc)}.VfPpkd-IkaYrd:hover .VfPpkd-Jh9lGc::before,.VfPpkd-IkaYrd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.VfPpkd-TolmDb{color:rgba(255,255,255,.87)}.VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgba(255,255,255,.87);background-color:var(--mdc-ripple-color,rgba(255,255,255,.87))}.VfPpkd-TolmDb:hover .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-TolmDb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{transition:opacity .15s linear}.VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.VfPpkd-TolmDb.VfPpkd-TolmDb{width:36px;height:36px;padding:6px;font-size:18px}.VfPpkd-TolmDb.VfPpkd-TolmDb .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:36px;max-width:36px}.VfPpkd-TolmDb.VfPpkd-TolmDb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:36px;height:36px;margin-top:0;margin-bottom:0;margin-right:0;margin-left:0}.VfPpkd-TolmDb.VfPpkd-TolmDb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:36px;max-width:36px}.VfPpkd-TolmDb.VfPpkd-TolmDb .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:36px;left:50%;width:36px;transform:translate(-50%,-50%)}.VOBzC{margin:24px}.VOBzC .VfPpkd-YAxtVc{background-color:rgb(32,33,36)}.VOBzC .VfPpkd-gIZMF{color:rgb(232,234,237)}.VOBzC .VfPpkd-IkaYrd:not(:disabled){background-color:transparent}.VOBzC .VfPpkd-IkaYrd:not(:disabled){color:rgb(138,180,248);color:var(--gm-colortextbutton-ink-color,rgb(138,180,248))}.VOBzC .VfPpkd-IkaYrd:disabled{color:rgba(232,234,237,.38);color:var(--gm-colortextbutton-disabled-ink-color,rgba(232,234,237,.38))}.VOBzC .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.VOBzC .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(138,180,248)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VOBzC .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.VOBzC .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.VOBzC .VfPpkd-IkaYrd:hover:not(:disabled),.VOBzC .VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.VOBzC .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.VOBzC .VfPpkd-IkaYrd:active:not(:disabled){color:rgb(174,203,250);color:var(--gm-colortextbutton-ink-color--stateful,rgb(174,203,250))}.VOBzC .VfPpkd-IkaYrd .VfPpkd-Jh9lGc::before,.VOBzC .VfPpkd-IkaYrd .VfPpkd-Jh9lGc::after{background-color:rgb(174,203,250);background-color:var(--gm-colortextbutton-state-color,rgb(174,203,250))}.VOBzC .VfPpkd-IkaYrd:hover .VfPpkd-Jh9lGc::before,.VOBzC .VfPpkd-IkaYrd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VOBzC .VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VOBzC .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VOBzC .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.VOBzC .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.VOBzC .VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.VOBzC .VfPpkd-TolmDb{color:rgb(232,234,237);z-index:0}.VOBzC .VfPpkd-TolmDb:hover .VfPpkd-Bz112c-Jh9lGc::before,.VOBzC .VfPpkd-TolmDb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.VOBzC .VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.VOBzC .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.VOBzC .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.VOBzC .VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.VOBzC .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::before,.VOBzC .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.VOBzC .VfPpkd-TolmDb:disabled{color:rgba(232,234,237,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(232,234,237,.38))}.VOBzC .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::before,.VOBzC .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.VOBzC .VfPpkd-TolmDb:hover .VfPpkd-Bz112c-Jh9lGc::before,.VOBzC .VfPpkd-TolmDb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VOBzC .VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.VOBzC .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VOBzC .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{transition:opacity .15s linear}.VOBzC .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.VOBzC .VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.VOBzC .VfPpkd-TolmDb{width:36px;height:36px;padding:6px}.VOBzC .VfPpkd-TolmDb .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:36px;max-width:36px}.VOBzC .VfPpkd-TolmDb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:36px;height:36px;margin-top:0;margin-bottom:0;margin-right:0;margin-left:0}.VOBzC .VfPpkd-TolmDb.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:36px;max-width:36px}.VOBzC .VfPpkd-TolmDb .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:36px;left:50%;width:36px;transform:translate(-50%,-50%)}.Uo6OHe{background:transparent;max-width:47.5rem;width:100%;overflow-y:auto}.Uo6OHe>[jsslot]{-moz-border-radius:0.5rem;border-radius:0.5rem}.mgGKnc{width:15.625rem}.NfDqfe{width:100%}.gWB1lc{width:100%}.GXzb2d{width:100%}.lsZcSc{margin:-0.5rem -1rem}.uRr8Jb .Fxmcue{padding:0.75rem;padding-left:1rem}.uRr8Jb .snByac{font-family:Roboto,Arial,sans-serif;font-size:14px;font-weight:400;letter-spacing:.2px;line-height:20px;margin-right:0.25rem}.uRr8Jb:not(.RDPZE) .snByac{color:#202124}.Kx1b0{height:1.5rem;margin-right:0.5rem;width:1.5rem}.SBgUnc{margin-bottom:1rem}.mNfPw{margin-top:1rem}.LJx7of{background-color:#f8f9fa}.LJx7of.enlinc .Fxmcue{align-items:center;box-sizing:border-box;display:-webkit-inline-box;display:-webkit-inline-flex;display:-ms-inline-flexbox;display:inline-flex;justify-content:space-between;text-align:left;width:100%}.Oz1VGd{color:#9aa0a6}.Z99Cif{word-break:break-all}.WGcIBc{margin-bottom:1rem}.Oh6Vl{margin-bottom:1rem;margin-top:1rem}.qOzNpe{margin-left:0.5rem;width:auto}.qOzNpe .EmVfjc{height:18px;width:18px}.FMIZ6c{justify-content:flex-end}.FMIZ6c>div{margin-left:1rem}.meyvr{border-top:0.0625rem solid #e0e0e0;margin:0 -1rem;padding:1rem}.m6f1N{width:100%}.UtFhj{margin-top:0.5rem}.klG8ee{margin-right:0.5rem}.HFYDF{-moz-flex-wrap:wrap;flex-wrap:wrap;margin-top:-1rem}.HFYDF>div{margin-top:1rem}.pdwdEb{margin-right:1rem}.SbnRSc.SbnRSc{-moz-box-sizing:border-box;box-sizing:border-box;max-height:100%;max-width:100%}.SbnRSc .wnIM7{-moz-box-sizing:border-box;box-sizing:border-box;height:34.375rem;max-height:100%;max-width:100%;padding:0;width:47.25rem}.TDg32e{height:100%}.sjgYwf{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;height:100%;overflow:hidden}.ISy4H{-moz-box-align:center;align-items:center;-moz-box-sizing:border-box;box-sizing:border-box;display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;-moz-box-flex:0;flex:0 0 auto;padding:1.5rem;width:100%}.iPtkNb{margin-right:1rem}.aHMLCc{display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;margin-top:-.5rem;padding:.5rem 1.5rem}.cmTiyd{border-top:.0625rem solid rgb(218,220,224);-moz-box-flex:1;flex:1 1 auto;overflow:auto}.t5tYqf .cmTiyd{border-bottom:.0625rem solid rgb(218,220,224)}.pGPH1e{padding:.5rem 1.5rem}.XDSyOc{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-flex:0;flex:0 0 auto;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;-moz-box-pack:justify;justify-content:space-between;padding:1.5rem}.T4pcrc{padding:.5rem 1.5rem}.pGPH1e .aGtBAd{width:100%}.pGPH1e .YfHqed{display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;width:100%}.XlStVe,.NzjwC,.PiOU2e{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;-moz-box-orient:horizontal;-moz-box-direction:normal;flex-direction:row;-moz-box-flex:0;flex-grow:0;flex-shrink:0;overflow:hidden;width:100%}.XlStVe{flex-basis:20.625rem;padding-right:1rem}.ErXmq{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;height:100%;margin-right:.75rem}.ErXmq .tkmmwb{align-self:center}.ARHFvd{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;overflow:hidden}.NzjwC{flex-basis:13.75rem;padding-right:1rem}.PiOU2e{flex-basis:6.875rem;margin-right:1rem}.FqHKUe.FqHKUe .dNuvt{padding:1rem}.NETtEe{display:none}@media (max-width:870px){.NETtEe{display:block}.aHMLCc{display:none}.pGPH1e{padding:.5rem 1rem}.XlStVe{flex-basis:100%}.NzjwC,.PiOU2e{display:none}}.gpeXDe{border-bottom:.0625rem solid rgb(218,220,224);margin:0 -1rem 1.5rem;padding:1rem}.lIZXM{margin-top:1rem;width:100%}.lIZXM:not(.mKfy1){flex-wrap:wrap}.i84rE,.U1rsQb{flex-shrink:0}.U1rsQb.oxacD{margin-left:0}.TPWgGb.TPWgGb{margin-right:-1rem}.azralf{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;margin-top:2rem}.rjGFOb{max-width:100%;width:47.5rem}.g37tgd{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.CSivxe{background-color:#f1f3f4;padding:2rem}.u9RzIb{margin-top:1rem;max-width:24.0625rem}.y7i1Nc{margin-bottom:1rem;width:6.25rem}.d2b4L{padding:1.5rem}.U71Lnc{margin-bottom:1.5rem}.VMWAxd{margin-top:2rem}.RInnx{text-align:center;width:100%}.L167uf{margin:0 0.5rem 0 1rem}.nbFnZ{margin:1rem 0}.ZbysJe{margin-bottom:1rem}.WEjkH.WEjkH{display:inline-block;margin-top:0}.dbsF4b .qRUolc{text-align:center}.dbsF4b .J9fJmf{flex-direction:row-reverse;justify-content:end}.L6Tcab{color:#d50000}.Ka95Z{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.EaTUdc,.UmX19b{margin-left:1rem;width:8.125rem}@media (max-width:30em){.oz51Ne{width:6.875rem}.EaTUdc,.UmX19b{width:5.625rem}}.Ka95Z .aCsJod.oJeWuf{padding-top:1rem}.EWKrtf{margin-top:1rem}.RxsGPe:empty{display:none}.yFza7b{height:52px}.DS3fne{color:rgb(154,160,166)}.apFhrb{margin-right:1rem;width:11.25rem}.suIOVe{-moz-box-align:start;align-items:flex-start;display:-moz-box;display:flex;flex-wrap:no-wrap;margin-bottom:1rem;padding-right:.125rem}.DqmUvd{margin-top:-0.25rem}.H1keZd{margin-bottom:1rem}.PfUTwd{color:#d50000}.Gmvs1{display:inline-block;margin-top:0.25rem;text-align:right;width:200px}.XUcbLe{display:inline-block;margin-left:1rem}.Gf7iTb:empty{margin-top:-1.5rem}.kzJRP{margin:0.5rem 0;margin-left:-0.5rem}.AHZqAf .vUBwW{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;color:#fff;height:2.5rem;line-height:2.5rem;margin-left:-.625rem;text-transform:uppercase;width:2.5rem}.DC43lf .vUBwW{margin-top:-1.5rem}.g6gble{-moz-box-align:center;align-items:center;display:-moz-box;display:flex;overflow:hidden}.QeGaRd{padding-bottom:.25rem;padding-top:.25rem}.jYRzx{padding-bottom:1rem}.wgdZlc{font-family:Roboto,Arial,sans-serif;line-height:1rem;font-size:.75rem;letter-spacing:.025em;font-weight:400;color:rgb(95,99,104);left:3.5rem;position:fixed}.pixFV{bottom:1.875rem;display:-moz-box;display:flex;padding:.3125rem;position:fixed}.zevhc{bottom:1.5rem;display:-moz-box;display:flex;padding:.3125rem;position:fixed}.FzFOE{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;color:rgb(60,64,67)}.I6N0E{max-height:33.4375rem;min-width:35.3125rem}@media (max-width:40rem){.I6N0E{min-width:29.0625rem}}@media (max-width:30rem){.I6N0E{min-width:23.75rem}}.pC9vb{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400;color:rgb(95,99,104)}.Lz37cd{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:500}.VfPpkd-Cv7pCf{position:relative;display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;width:328px;overflow:hidden}.VfPpkd-npdOxb{z-index:9000}.VfPpkd-Cv7pCf-tJHJj{display:-moz-box;display:flex;-moz-box-pack:justify;justify-content:space-between;padding:8px}.VfPpkd-UrYcU-XnnMxf-EglORb{position:absolute;top:-9999px;left:-9999px;height:1px;overflow:hidden;font-size:0}.VfPpkd-HhDot-tJHJj-eEDwDf{padding:0}.VfPpkd-HhDot-tJHJj{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit);width:44px;height:44px;line-height:44px}.VfPpkd-XqMb-JNdkSc{display:-moz-box;display:flex;-moz-box-pack:justify;justify-content:space-between}.VfPpkd-XqMb-hFsbo{width:44px;height:44px;padding:10px;margin:2px 0}.VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:44px;max-width:44px}.VfPpkd-XqMb-hFsbo.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:40px;height:40px;margin-top:2px;margin-bottom:2px;margin-right:2px;margin-left:2px}.VfPpkd-XqMb-hFsbo.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:40px;max-width:40px}.VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:44px;left:50%;width:44px;transform:translate(-50%,-50%)}.VfPpkd-XqMb-S2QgGf-kj0dLd{padding-left:4px;padding-right:0;min-width:0}[dir=rtl] .VfPpkd-XqMb-S2QgGf-kj0dLd,.VfPpkd-XqMb-S2QgGf-kj0dLd[dir=rtl]{padding-left:0;padding-right:4px}.VfPpkd-XqMb-S2QgGf-kj0dLd .VfPpkd-kBDsod{margin:0;width:24px;height:24px}.VfPpkd-XqMb-S2QgGf-kj0dLd:disabled .VfPpkd-kBDsod{visibility:hidden}.VfPpkd-XqMb-hFsbo,.VfPpkd-XqMb-S2QgGf-kj0dLd{z-index:1}.VfPpkd-hOoMI-haAclf{visibility:hidden;height:calc(100% - 8px);width:100%;position:absolute;top:0;overflow:auto}.VfPpkd-hOoMI{position:relative;-moz-box-sizing:border-box;box-sizing:border-box;min-height:100%}.VfPpkd-hOoMI-ibnC6b .VfPpkd-rymPhb-pZXsl::before{opacity:0}.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:40px}.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:48px}.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:64px}.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b,.VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-hOoMI-ibnC6b .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-hOoMI-ibnC6b .VfPpkd-rymPhb-KkROqb,.VfPpkd-hOoMI-ibnC6b .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf,.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf{border-top:1px solid}.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-Cv7pCf-jyrRxf,.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-Cv7pCf-qJTHM,.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-Cv7pCf-jyrRxf,.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-Cv7pCf-qJTHM{visibility:hidden}.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf,.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf{visibility:visible}.VfPpkd-hOoMI-ibnC6b-barxie-Bz112c{visibility:hidden}.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-hOoMI-ibnC6b-barxie-Bz112c{visibility:visible}.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-XqMb-hFsbo,.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-XqMb-hFsbo{visibility:hidden}.VfPpkd-Cv7pCf-qJTHM{position:relative}.VfPpkd-Cv7pCf-jyrRxf{margin:0 10px 4px;width:calc(100% - 20px);border-spacing:0}.VfPpkd-BE01ge-eEDwDf{width:44px;height:44px}.VfPpkd-RKhZBe-eEDwDf{padding:0}.VfPpkd-RKhZBe-LgbsSe{width:36px;height:36px;min-width:0;padding:0;border:none;border-radius:18px;margin-top:4px;margin-bottom:4px;margin-right:4px;margin-left:4px}.VfPpkd-RKhZBe-LgbsSe.VfPpkd-RKhZBe-LgbsSe.VfPpkd-LgbsSe{font-family:var(--mdc-typography-font-family,Roboto,sans-serif);-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-moz-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit);font-weight:500;font-size:.75rem}.VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc{border-radius:18px}.VfPpkd-RKhZBe-LgbsSe .VfPpkd-RLmnJb{position:absolute;top:50%;height:44px;left:50%;width:44px;transform:translate(-50%,-50%)}.VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:hover{cursor:default}.VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe.VfPpkd-LgbsSe,.VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me.VfPpkd-RKhZBe-LgbsSe.VfPpkd-LgbsSe,.VfPpkd-RKhZBe-LgbsSe:disabled.VfPpkd-RKhZBe-LgbsSe.VfPpkd-LgbsSe{font-weight:400}.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l{border:1px solid}.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd{border:none}.VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::after{top:0;left:0;width:100%;height:100%}.VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc.VfPpkd-ksKsZd-mWPk3d::before,.VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc.VfPpkd-ksKsZd-mWPk3d::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0);width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc.VfPpkd-ksKsZd-mWPk3d::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-RKhZBe-eEDwDf .VfPpkd-dgl2Hf-ppHlrf-sM5MNb{pointer-events:none;position:relative;z-index:0}.VfPpkd-RKhZBe-LgbsSe{will-change:unset;pointer-events:auto}.VfPpkd-RKhZBe-LgbsSe .VfPpkd-RLmnJb{z-index:-1}.VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc{pointer-events:none}.VfPpkd-Cv7pCf-LQLjdd{display:-moz-box;display:flex;height:52px}.VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus{outline:1px solid transparent}@media screen and (forced-colors:active){.VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus{outline-color:CanvasText}}.VfPpkd-XqMb-hFsbo.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-XqMb-hFsbo:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-XqMb-hFsbo.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-XqMb-hFsbo:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{border-color:CanvasText}}.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:3px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd::before{border-color:CanvasText}}.VfPpkd-XqMb-S2QgGf-kj0dLd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-XqMb-S2QgGf-kj0dLd:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-XqMb-S2QgGf-kj0dLd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-XqMb-S2QgGf-kj0dLd:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{border-color:CanvasText}}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me,.VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me{color:GrayText}}@media (max-width:328px){.VfPpkd-Cv7pCf{width:320px}.VfPpkd-Cv7pCf-tJHJj{padding:8px 4px}.VfPpkd-Cv7pCf-jyrRxf{margin:0 6px 4px;width:calc(100% - 12px)}}.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-Jh9lGc::after{background-color:#000;background-color:var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me{color:rgba(0,0,0,.38)}.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:hover,.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:not(.VfPpkd-ksKsZd-mWPk3d):focus,.VfPpkd-Cv7pCf .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:not(:disabled):active{color:rgba(0,0,0,.38)}.VfPpkd-Cv7pCf .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){color:#000;color:var(--mdc-text-button-label-text-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-XqMb-S2QgGf-kj0dLd:disabled{color:#000;color:var(--mdc-text-button-disabled-label-text-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:transparent}.VfPpkd-Cv7pCf .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.VfPpkd-Cv7pCf .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-hOoMI-haAclf{background-color:white}.VfPpkd-Cv7pCf.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled),.VfPpkd-Cv7pCf.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){color:#000;color:var(--mdc-text-button-label-text-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled),.VfPpkd-Cv7pCf.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){background-color:rgba(0,0,0,.12)}.VfPpkd-Cv7pCf.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf,.VfPpkd-Cv7pCf.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf{border-top-color:#bdbdbd}.VfPpkd-Cv7pCf .VfPpkd-HhDot-tJHJj{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe:not(:disabled){color:#000;color:var(--mdc-outlined-button-label-text-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe:disabled{color:rgba(0,0,0,.38);color:var(--mdc-outlined-button-disabled-label-text-color,rgba(0,0,0,.38))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::after{background-color:#000;background-color:var(--mdc-outlined-button-hover-state-layer-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){color:#6200ee;color:var(--mdc-outlined-button-label-text-color,var(--mdc-theme-primary,#6200ee))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::before,.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::after{background-color:#6200ee;background-color:var(--mdc-outlined-button-hover-state-layer-color,var(--mdc-theme-primary,#6200ee))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){border-color:#6200ee;border-color:var(--mdc-outlined-button-outline-color,var(--mdc-theme-primary,#6200ee))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){color:#fff;color:var(--mdc-outlined-button-label-text-color,var(--mdc-theme-surface,#fff))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::before,.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::after{background-color:#000;background-color:var(--mdc-outlined-button-hover-state-layer-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){background-color:#6200ee;background-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled){color:rgba(0,0,0,.38);color:var(--mdc-outlined-button-label-text-color,rgba(0,0,0,.38))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):hover{color:rgba(0,0,0,.38);color:var(--mdc-outlined-button-hover-label-text-color,rgba(0,0,0,.38))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgba(0,0,0,.38);color:var(--mdc-outlined-button-focus-label-text-color,rgba(0,0,0,.38))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):not(:disabled):active{color:rgba(0,0,0,.38);color:var(--mdc-outlined-button-pressed-label-text-color,rgba(0,0,0,.38))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled){color:rgba(0,0,0,.38);color:var(--mdc-outlined-button-label-text-color,rgba(0,0,0,.38))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){color:#6200ee;color:var(--mdc-outlined-button-label-text-color,var(--mdc-theme-primary,#6200ee))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::before,.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::after{background-color:#6200ee;background-color:var(--mdc-outlined-button-hover-state-layer-color,var(--mdc-theme-primary,#6200ee))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){border-color:#6200ee;border-color:var(--mdc-outlined-button-outline-color,var(--mdc-theme-primary,#6200ee))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){color:#fff;color:var(--mdc-outlined-button-label-text-color,var(--mdc-theme-surface,#fff))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::before,.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::after{background-color:#000;background-color:var(--mdc-outlined-button-hover-state-layer-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Cv7pCf .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){background-color:#6200ee;background-color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-t0sizb{border-radius:8px;max-width:none;max-height:none}.VfPpkd-t0sizb .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-t0sizb::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-t0sizb::before{border-color:CanvasText}}.VfPpkd-PFym2e-LgbsSe-haAclf,.VfPpkd-eSiNeb-JIbuQc{margin-left:16px;margin-right:0}[dir=rtl] .VfPpkd-PFym2e-LgbsSe-haAclf,[dir=rtl] .VfPpkd-eSiNeb-JIbuQc,.VfPpkd-PFym2e-LgbsSe-haAclf[dir=rtl],.VfPpkd-eSiNeb-JIbuQc[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-eSiNeb-IbE0S-LgbsSe-haAclf{margin-left:auto;margin-right:16px}[dir=rtl] .VfPpkd-eSiNeb-IbE0S-LgbsSe-haAclf,.VfPpkd-eSiNeb-IbE0S-LgbsSe-haAclf[dir=rtl]{margin-left:16px;margin-right:auto}.VfPpkd-GRS59e{min-width:44px}.VfPpkd-GRS59e.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{position:absolute;-moz-box-sizing:border-box;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-GRS59e.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{border-color:CanvasText}}@media (max-width:328px){.VfPpkd-PFym2e-LgbsSe-haAclf,.VfPpkd-eSiNeb-JIbuQc{margin-left:12px;margin-right:0}[dir=rtl] .VfPpkd-PFym2e-LgbsSe-haAclf,[dir=rtl] .VfPpkd-eSiNeb-JIbuQc,.VfPpkd-PFym2e-LgbsSe-haAclf[dir=rtl],.VfPpkd-eSiNeb-JIbuQc[dir=rtl]{margin-left:0;margin-right:12px}.VfPpkd-eSiNeb-IbE0S-LgbsSe-haAclf{margin-left:auto;margin-right:12px}[dir=rtl] .VfPpkd-eSiNeb-IbE0S-LgbsSe-haAclf,.VfPpkd-eSiNeb-IbE0S-LgbsSe-haAclf[dir=rtl]{margin-left:12px;margin-right:auto}}.VfPpkd-t0sizb .VfPpkd-GRS59e:not(:disabled){color:#6200ee;color:var(--mdc-text-button-label-text-color,var(--mdc-theme-primary,#6200ee))}.VfPpkd-t0sizb .VfPpkd-GRS59e .VfPpkd-Jh9lGc::before,.VfPpkd-t0sizb .VfPpkd-GRS59e .VfPpkd-Jh9lGc::after{background-color:#6200ee;background-color:var(--mdc-text-button-hover-state-layer-color,var(--mdc-theme-primary,#6200ee))}.bc5ALd .VfPpkd-XqMb-hFsbo{color:rgb(95,99,104)}.bc5ALd .VfPpkd-XqMb-hFsbo:hover{color:rgb(32,33,36)}.bc5ALd .VfPpkd-XqMb-hFsbo.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-XqMb-hFsbo:not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36)}.bc5ALd .VfPpkd-XqMb-hFsbo:not(:disabled):active{color:rgb(32,33,36)}.bc5ALd .VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-Jh9lGc::before,.bc5ALd .VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.bc5ALd .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me{color:rgba(60,64,67,.38)}.bc5ALd .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:hover,.bc5ALd .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:not(.VfPpkd-ksKsZd-mWPk3d):focus,.bc5ALd .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:not(:disabled):active{color:rgba(60,64,67,.38)}.bc5ALd .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){color:rgb(95,99,104);color:var(--mdc-text-button-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled):hover{color:rgb(32,33,36);color:var(--mdc-text-button-hover-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36);color:var(--mdc-text-button-focus-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled):not(:disabled):active{color:rgb(32,33,36);color:var(--mdc-text-button-pressed-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-XqMb-S2QgGf-kj0dLd:disabled{color:rgb(95,99,104);color:var(--mdc-text-button-disabled-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:transparent}.bc5ALd .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.bc5ALd .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.bc5ALd .VfPpkd-hOoMI-haAclf{background-color:#fff}.bc5ALd.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled),.bc5ALd.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){color:rgb(32,33,36);color:var(--mdc-text-button-label-text-color,rgb(32,33,36))}.bc5ALd.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled),.bc5ALd.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){background-color:rgba(60,64,67,.12)}.bc5ALd.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf,.bc5ALd.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf{border-top-color:rgb(218,220,224)}.bc5ALd .VfPpkd-HhDot-tJHJj{color:rgb(95,99,104)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(:disabled){color:rgb(60,64,67);color:var(--mdc-outlined-button-label-text-color,rgb(60,64,67))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(:disabled):hover{color:rgb(32,33,36);color:var(--mdc-outlined-button-hover-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36);color:var(--mdc-outlined-button-focus-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(:disabled):not(:disabled):active{color:rgb(32,33,36);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:disabled{color:rgb(95,99,104);color:var(--mdc-outlined-button-disabled-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::after{background-color:rgb(60,64,67);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(60,64,67))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:hover .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.04)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.12)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.bc5ALd .VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.1)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.1)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){color:rgb(26,115,232);color:var(--mdc-outlined-button-label-text-color,rgb(26,115,232))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{color:rgb(23,78,166);color:var(--mdc-outlined-button-hover-label-text-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(23,78,166);color:var(--mdc-outlined-button-focus-label-text-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(:disabled):active{color:rgb(23,78,166);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::after{background-color:rgb(23,78,166);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:hover .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.04)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.12)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.1)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.1)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){border-color:rgb(26,115,232);border-color:var(--mdc-outlined-button-outline-color,rgb(26,115,232))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(23,78,166);border-color:var(--mdc-outlined-button-focus-outline-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{border-color:rgb(23,78,166)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):active,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):focus:active{border-color:rgb(23,78,166)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){color:#fff;color:var(--mdc-outlined-button-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{color:#fff;color:var(--mdc-outlined-button-hover-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:#fff;color:var(--mdc-outlined-button-focus-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{color:#fff;color:var(--mdc-outlined-button-pressed-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:hover .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.16;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.16)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.24)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.2;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.2)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.2)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){background-color:rgb(26,115,232)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{background-color:rgb(26,115,232)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{background-color:rgb(26,115,232)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{background-color:rgb(26,115,232)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled){color:rgb(95,99,104);color:var(--mdc-outlined-button-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):hover{color:rgb(95,99,104);color:var(--mdc-outlined-button-hover-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(95,99,104);color:var(--mdc-outlined-button-focus-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):not(:disabled):active{color:rgb(95,99,104);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled){color:rgb(95,99,104);color:var(--mdc-outlined-button-label-text-color,rgb(95,99,104))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled):hover{color:rgb(32,33,36);color:var(--mdc-outlined-button-hover-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36);color:var(--mdc-outlined-button-focus-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled):not(:disabled):active{color:rgb(32,33,36);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){color:rgb(26,115,232);color:var(--mdc-outlined-button-label-text-color,rgb(26,115,232))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{color:rgb(23,78,166);color:var(--mdc-outlined-button-hover-label-text-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(23,78,166);color:var(--mdc-outlined-button-focus-label-text-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(:disabled):active{color:rgb(23,78,166);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::after{background-color:rgb(23,78,166);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:hover .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.04)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.12)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.1)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.1)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){border-color:rgb(26,115,232);border-color:var(--mdc-outlined-button-outline-color,rgb(26,115,232))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(23,78,166);border-color:var(--mdc-outlined-button-focus-outline-color,rgb(23,78,166))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{border-color:rgb(23,78,166)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):active,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):focus:active{border-color:rgb(23,78,166)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){color:#fff;color:var(--mdc-outlined-button-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{color:#fff;color:var(--mdc-outlined-button-hover-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:#fff;color:var(--mdc-outlined-button-focus-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{color:#fff;color:var(--mdc-outlined-button-pressed-label-text-color,#fff)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(32,33,36))}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:hover .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.16;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.16)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.24;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.24)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.2;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.2)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.2)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){background-color:rgb(26,115,232)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{background-color:rgb(26,115,232)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{background-color:rgb(26,115,232)}.bc5ALd .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{background-color:rgb(26,115,232)}.uIJlfe{z-index:2051}.uIJlfe .VfPpkd-GRS59e:not(:disabled){color:rgb(26,115,232);color:var(--mdc-text-button-label-text-color,rgb(26,115,232))}.uIJlfe .VfPpkd-GRS59e:not(:disabled):hover{color:rgb(23,78,166);color:var(--mdc-text-button-hover-label-text-color,rgb(23,78,166))}.uIJlfe .VfPpkd-GRS59e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.uIJlfe .VfPpkd-GRS59e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(23,78,166);color:var(--mdc-text-button-focus-label-text-color,rgb(23,78,166))}.uIJlfe .VfPpkd-GRS59e:not(:disabled):not(:disabled):active{color:rgb(23,78,166);color:var(--mdc-text-button-pressed-label-text-color,rgb(23,78,166))}.uIJlfe .VfPpkd-GRS59e .VfPpkd-Jh9lGc::before,.uIJlfe .VfPpkd-GRS59e .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--mdc-text-button-hover-state-layer-color,rgb(26,115,232))}.uIJlfe .VfPpkd-GRS59e:hover .VfPpkd-Jh9lGc::before,.uIJlfe .VfPpkd-GRS59e.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-text-button-hover-state-layer-opacity,.04)}.uIJlfe .VfPpkd-GRS59e.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.uIJlfe .VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{transition-duration:75ms;opacity:.12;opacity:var(--mdc-text-button-focus-state-layer-opacity,.12)}.uIJlfe .VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{transition:opacity .15s linear}.uIJlfe .VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{transition-duration:75ms;opacity:.1;opacity:var(--mdc-text-button-pressed-state-layer-opacity,.1)}.uIJlfe .VfPpkd-GRS59e.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-text-button-pressed-state-layer-opacity,0.1)}.VfPpkd-Zc28rc{display:-moz-inline-box;display:inline-flex;position:relative}.VfPpkd-Zc28rc[hidden]{display:none}.VfPpkd-Cv7pCf-ornU0b{border-radius:50%;transition:75ms background-color linear}.VfPpkd-Cv7pCf-ornU0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-Cv7pCf-ornU0b:not(.VfPpkd-ksKsZd-mWPk3d):focus{outline:1px solid transparent}@media screen and (forced-colors:active){.VfPpkd-Cv7pCf-ornU0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-Cv7pCf-ornU0b:not(.VfPpkd-ksKsZd-mWPk3d):focus{outline-color:CanvasText}}.VfPpkd-Cv7pCf-ornU0b-sM5MNb{position:absolute;top:6px;left:auto;right:0}[dir=rtl] .VfPpkd-Cv7pCf-ornU0b-sM5MNb,.VfPpkd-Cv7pCf-ornU0b-sM5MNb[dir=rtl]{left:0;right:auto}.VfPpkd-oEZKA-H9tDt,.VfPpkd-Ugjwi{width:100%}.VfPpkd-oEZKA-YPqjbf{margin-left:0;margin-right:56px}[dir=rtl] .VfPpkd-oEZKA-YPqjbf,.VfPpkd-oEZKA-YPqjbf[dir=rtl]{margin-left:56px;margin-right:0}.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b:hover .VfPpkd-Bz112c-Jh9lGc::before{opacity:.12}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-oEZKA{height:56px}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b-sM5MNb{margin:0 6px;max-width:44px;max-height:44px}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b{width:44px;height:44px;padding:10px}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:44px;max-width:44px}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:40px;height:40px;margin-top:2px;margin-bottom:2px;margin-right:2px;margin-left:2px}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:40px;max-width:40px}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:44px;left:50%;width:44px;transform:translate(-50%,-50%)}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(0,0,0,.38)}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::after{background-color:#000;background-color:var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Zc28rc-OWXEXe-MFS4be.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b{background-color:rgba(0,0,0,.12)}.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-Cv7pCf-ornU0b:hover:disabled,.VfPpkd-Zc28rc-OWXEXe-MFS4be .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(0,0,0,.38)}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA{height:56px}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-37.25px) scale(1)}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:.75rem}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{transform:translateY(-34.75px) scale(.75)}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA.VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe,.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA .VfPpkd-NSFCdd-i5vt6e-OWXEXe-mWPk3d .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{font-size:1rem}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA .VfPpkd-NLUYnc-V67aGc-OWXEXe-bF1zU{animation:mdc-floating-label-shake-float-above-text-field-outlined-56px .25s 1}@keyframes mdc-floating-label-shake-float-above-text-field-outlined-56px{0%{transform:translateX(0) translateY(-34.75px) scale(.75)}33%{animation-timing-function:cubic-bezier(.5,0,.701732,.495819);transform:translateX(4%) translateY(-34.75px) scale(.75)}66%{animation-timing-function:cubic-bezier(.302435,.381352,.55,.956352);transform:translateX(-4%) translateY(-34.75px) scale(.75)}100%{transform:translateX(0) translateY(-34.75px) scale(.75)}}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b-sM5MNb{margin:0 6px;max-width:44px;max-height:44px}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b{width:44px;height:44px;padding:10px}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:44px;max-width:44px}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:40px;height:40px;margin-top:2px;margin-bottom:2px;margin-right:2px;margin-left:2px}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:40px;max-width:40px}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:44px;left:50%;width:44px;transform:translate(-50%,-50%)}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(0,0,0,.38)}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::after{background-color:#000;background-color:var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Zc28rc-OWXEXe-INsAgc.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b{background-color:rgba(0,0,0,.12)}.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-Cv7pCf-ornU0b:hover:disabled,.VfPpkd-Zc28rc-OWXEXe-INsAgc .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(0,0,0,.38)}.a0QCRb .VfPpkd-Cv7pCf-ornU0b{color:rgb(95,99,104)}.a0QCRb .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(95,99,104,.38)}.a0QCRb .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::before,.a0QCRb .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.a0QCRb .VfPpkd-Cv7pCf-ornU0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.a0QCRb .VfPpkd-Cv7pCf-ornU0b:not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36)}.a0QCRb .VfPpkd-Cv7pCf-ornU0b:not(:disabled):active{color:rgb(32,33,36)}.a0QCRb.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b{color:rgb(32,33,36);background-color:rgba(60,64,67,.12)}.a0QCRb .VfPpkd-Cv7pCf-ornU0b:hover,.a0QCRb .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b{color:rgb(32,33,36)}.a0QCRb .VfPpkd-Cv7pCf-ornU0b:hover:disabled,.a0QCRb .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(95,99,104,.38)}.xesam .VfPpkd-Cv7pCf-ornU0b{color:rgb(95,99,104)}.xesam .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(95,99,104,.38)}.xesam .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::before,.xesam .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.xesam .VfPpkd-Cv7pCf-ornU0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.xesam .VfPpkd-Cv7pCf-ornU0b:not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36)}.xesam .VfPpkd-Cv7pCf-ornU0b:not(:disabled):active{color:rgb(32,33,36)}.xesam.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b{color:rgb(32,33,36);background-color:rgba(60,64,67,.12)}.xesam .VfPpkd-Cv7pCf-ornU0b:hover,.xesam .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b{color:rgb(32,33,36)}.xesam .VfPpkd-Cv7pCf-ornU0b:hover:disabled,.xesam .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(95,99,104,.38)}.RZ2Y3.oJ9Ind .VfPpkd-oEZKA{height:52px}.RZ2Y3.oJ9Ind .VfPpkd-Cv7pCf-ornU0b-sM5MNb{margin:0 8px;max-width:40px;max-height:40px}.RZ2Y3.oJ9Ind .VfPpkd-Cv7pCf-ornU0b{width:40px;height:40px;padding:8px}.RZ2Y3.oJ9Ind .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:40px;max-width:40px}.RZ2Y3.oJ9Ind .VfPpkd-Cv7pCf-ornU0b.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:40px;height:40px;margin-top:0;margin-bottom:0;margin-right:0;margin-left:0}.RZ2Y3.oJ9Ind .VfPpkd-Cv7pCf-ornU0b.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:40px;max-width:40px}.RZ2Y3.oJ9Ind .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:40px;left:50%;width:40px;transform:translate(-50%,-50%)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc,.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc,.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me).VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(197,34,31)}.mExmDc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(197,34,31)}.PIi4Cf{display:-moz-box;display:flex}@media (max-width:33.125rem){.PIi4Cf{display:inline-block}}.pkpPZc{color:rgb(154,160,166)}.oHIug{color:rgb(197,34,31)}.jTAjWd{-moz-box-align:start;align-items:flex-start;display:-moz-box;display:flex;flex-wrap:no-wrap;margin-top:1rem;padding-right:.125rem}.ptPUjc,.vpcS2b{margin-right:1rem;width:11.25rem}@media (max-width:33.125rem){.ptPUjc{width:15.625rem}}@media (max-width:50rem){.vpcS2b{width:23.5rem}}@media (max-width:33.125rem){.vpcS2b{width:15rem}}.oxBPSd{display:-moz-box;display:flex}@media (max-width:50rem){.oxBPSd{display:inline-block;padding-bottom:.5rem}}.ebLi5c{height:52px}.xLjkBc{flex-shrink:0}.hHxPyf{width:10rem}.rIRHO{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;color:rgb(60,64,67)}.js7GQd{margin-bottom:1rem;margin-top:1rem}.RPPiPc{margin-left:-.5rem}.tmY6ac{margin-bottom:1rem}.OKbzo{display:none;left:0;position:fixed;right:0;top:3.5rem}.ckIUie .OKbzo{display:block}.uR9cVd.oJeWuf{padding:0}.SHwQZd{margin:0 auto;max-width:700px;padding:1.5rem}@media (max-width:30em){.SHwQZd{padding:0.5rem}}.hwuvid{font-size:0.8125rem;margin-bottom:-1.5rem}@media (max-width:30em){.hwuvid{margin-bottom:-0.5rem}}.h50NT{line-height:0}.XKbOjc{padding:1.5rem;padding-bottom:0.5rem}.vO4eoc{margin-bottom:1.5rem}.SAKWs{margin-bottom:1rem}.vO4eoc~.vO4eoc,.SAKWs~.SAKWs{margin-top:2rem}.vO4eoc+.SAKWs{margin-top:0}.LqHDgc{border-bottom:0.0625rem solid #e0e0e0;margin:1.5rem -1rem 2rem}.cAO5X{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-flex-wrap:no-wrap;flex-wrap:no-wrap}.GeH8J{letter-spacing:.025em;font-family:Roboto,Arial,sans-serif;font-size:.75rem;font-weight:400;-moz-border-radius:3.25rem;border-radius:3.25rem;color:white;line-height:1.5rem;margin-left:0.5rem;margin-top:0.125rem;min-width:1.5rem;padding:0 0.375rem}.LjNQse{overflow:visible}.LjNQse .cTiNYb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-bottom:1rem}.LjNQse .tWfTvb{position:relative}.zt4tfb{margin-bottom:1.5rem}@charset "UTF-8";.tLBshf{width:20rem}.tLBshf .VfPpkd-TkwUic{height:40px;display:-moz-box;display:flex;-moz-box-align:baseline;align-items:baseline}.tLBshf .VfPpkd-TkwUic::before{display:inline-block;width:0;height:40px;content:"";vertical-align:0}.tLBshf .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS::before{content:"​"}.tLBshf .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS-haAclf{height:100%;display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center}.tLBshf .VfPpkd-TkwUic::before{display:none}.tLBshf .VfPpkd-TkwUic .VfPpkd-NLUYnc-V67aGc{display:none}.tLBshf.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS::before{content:"​"}.tLBshf.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic .VfPpkd-uusGie-fmcmS-haAclf{height:100%;display:-moz-inline-box;display:inline-flex;-moz-box-align:center;align-items:center}.tLBshf.VfPpkd-O1htCb-OWXEXe-di8rgd-V67aGc .VfPpkd-TkwUic::before{display:none}.tLBshf .VfPpkd-t08AT-Bz112c{width:20px;height:20px}.tLBshf.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc{max-width:calc(100% - 60px)}.tLBshf.VfPpkd-O1htCb-OWXEXe-MFS4be .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{max-width:calc(133.3333333333% - 80px)}.tLBshf .VfPpkd-StrnGf-rymPhb-ibnC6b,.tLBshf .VfPpkd-aJasdd-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:32px}.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:48px}.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-Gtdoyb{display:-moz-box;display:flex;-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column;-moz-box-pack:center;justify-content:center}.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS{margin-top:0;margin-bottom:0;line-height:1.4}.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS::before,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS::after{display:none}.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb,.tLBshf .VfPpkd-hjZysc-RWgCYc-wQNmvb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:56px}.WA09cf{margin:0.125rem 0}.hTD5hc{flex-shrink:0}.hKzOt{margin-bottom:1.5rem}@media (max-width:30rem){.hKzOt{display:block}}.PMLhsf:not(:empty){margin-top:0.5rem}.kzGuge{align-items:flex-start;padding:0.25rem 0.5rem}.IsRHDd{color:#a50e0e;margin-left:3rem}.ag5xxc{margin-left:3rem}.QPCpnf{align-items:center;color:#a50e0e;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;fill:#a50e0e;flex-shrink:0;padding-left:1.0625rem;width:1.4375rem}.gWxIGc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;gap:0.25rem;margin-top:0.125rem;width:19.75rem}@media (max-width:40em){.gWxIGc{width:15.625rem}}.GOGY4{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-flow:row wrap}.wlu0Lc{text-overflow:ellipsis;overflow:hidden;white-space:nowrap}.q8UhSb{padding-left:2.5rem}.G6I9Mb{text-align:right;width:3.25rem}.YdxQxe .wlu0Lc,.YdxQxe .G6I9Mb,.YdxQxe .vo2Wsc{color:#a50e0e}.OjzVP{margin-left:1rem;margin-top:0.25rem}.Tz6sTd{background-color:#f8f9fa;-moz-border-radius:0.5rem;border-radius:0.5rem;margin-bottom:0;margin-top:0.5rem}.Tz6sTd:first-of-type{margin-top:1rem}.Tz6sTd .JYB4b{padding:0.5rem 1rem}.PMLhsf .Tz6sTd[aria-expanded="true"] .JYB4b{border-bottom:0.0625rem solid #e0e0e0;margin-bottom:0.5rem}.lnpGb{margin:0 auto;max-width:43.75rem}.q4KgCc{left:0;position:fixed;right:0;top:3.5rem}.zo1Bhe{margin:0 0 1rem 1.5rem}.zo1Bhe .YrFhrf{margin-bottom:0.25rem}.ZvHxue{margin-bottom:0.5rem}.ZvHxue .JYB4b{color:#fff;background-color:#3c4043}.ZvHxue .D43mj{width:1.125rem}.ZvHxue .rKc6P{color:#fff;fill:#fff}.xVsAIc{padding:0.5rem 0}.xVsAIc ul{list-style:initial;margin:0.5rem 0;padding-left:2rem}.xVsAIc li{margin:0.5rem 0}.t0qXob{padding:1rem 1.5rem}.t0qXob:not(:last-of-type){border-bottom:0.0625rem solid #e0e0e0}.BDqqAe{background-color:#9aa0a6;height:2.25rem;margin-right:0.75rem;width:2.25rem}@media (max-width:40em){.uX0eBc{width:15.625rem}}.t0qXob.I8lGUd .BDqqAe{background-color:#a50e0e}.t0qXob.I8lGUd .LLP8tb{color:#a50e0e}.K4mNg{width:20rem}.Gjpklc{margin:0 0.25rem}.Gjpklc:last-of-type{display:none}.mxUcEe{margin-left:1.5rem}.owb53b{flex-direction:column}.xXsMpe{margin-bottom:0.5rem}.CyzZPb,.lVdIK{margin-bottom:1rem}.C7wCwf{list-style:disc;padding-left:1rem}.C7wCwf li:not(:last-child){margin-bottom:1rem}.xXsMpe{width:1.875rem}.S7nE7c{max-width:100%;width:448px}.O974kc{-moz-box-orient:vertical;-moz-box-direction:normal;flex-direction:column}.vxJi1c{display:block;margin:1rem auto 1.5rem;max-width:100%}.rw7Rv{margin-bottom:1rem}.lLZRtb{max-width:100%;width:50rem}.FVEPee{border-radius:.25rem;width:100%}.Nv6nWb{gap:1rem;flex-wrap:wrap;-moz-box-pack:justify;justify-content:space-between;margin-top:1.5rem}.ygw9c{flex-wrap:wrap;gap:1rem}.dH2B3c{margin-top:2rem}.jtUlhf{display:-moz-box;display:flex;flex-wrap:wrap;gap:.5rem;-moz-box-pack:justify;justify-content:space-between;margin-top:.5rem}.BRCGFd{border-radius:50%}.lHagT{color:#fff;fill:#fff}.BRCGFd[aria-checked=false] .lHagT{display:none}@media not all and (max-width:45em){.BRCGFd{height:4rem;width:4rem}.lHagT.lHagT{height:2rem;width:2rem}}sentinel{}</style><script async="" src="dec2_to_4_files/lazy.min.js" nonce=""></script><style nonce="" type="text/css" data-late-css="">.ZKQanf{margin-left:-0.25rem}sentinel{}</style><style nonce="" type="text/css" data-late-css="">.yJIkGf{padding:1rem 2rem}.pJFqib{display:-moz-box;display:flex;-moz-box-pack:center;justify-content:center;margin-bottom:2rem}.qa7ZLd{max-width:75%}.OcSfFd{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.5rem;font-weight:400;line-height:2rem}.ysWCZc{letter-spacing:.0142857143em;font-family:Roboto,Arial,sans-serif;font-size:.875rem;font-weight:400;line-height:1.25rem;padding:1rem 0}.pGryWb{margin-right:1rem}sentinel{}</style><style nonce="" type="text/css" data-late-css="">.mjbEJf{padding:1.5rem}.WLKmQe{margin-bottom:1rem}.SHkk9d{justify-content:flex-end}.SHkk9d>div{margin-left:1rem}sentinel{}</style><style nonce="" type="text/css" data-late-css="">.EbDdLe{font-style:italic;margin-top:.5rem}.wrkhkd{max-width:35rem}.be6XEc{margin-top:1rem}.Ae97qf{border:0;height:100%;width:100%}.yb5d6c{background:white;border-radius:8px;box-shadow:0 4px 16px rgba(0,0,0,.3);color:black;height:80%;outline:1px solid transparent;overflow:hidden;padding:0;position:fixed;width:80%;z-index:10001}@media (device-width:1024px) and (device-height:1366px) and (orientation:portrait),(device-width:1536px) and (device-height:2048px) and (orientation:portrait),(device-width:768px) and (device-height:1024px) and (orientation:portrait),(device-width:800px) and (device-height:1280px) and (orientation:portrait),(device-width:834px) and (device-height:1112px) and (orientation:portrait){.yb5d6c{height:45%;width:90%}}@media (max-device-height:480px),(max-device-width:640px){.yb5d6c{border-radius:0;height:100%;width:100%}}.yb5d6c-xJ5Hnf{background:#666;left:0;position:fixed;top:0;z-index:10000}.yb5d6c-bN97Pc{height:100%;width:100%}.yb5d6c-r4nke,.yb5d6c-r4nke-TvD9Pc{display:none}.BdlyXe{height:100%;width:100%;border-radius:0;transition:all .3s}sentinel{}</style><style nonce="" type="text/css" data-late-css="">.RM9ulf{visibility:hidden;position:fixed;z-index:5000;color:#fff;pointer-events:none}.RM9ulf.catR2e{max-width:90%;max-height:90%}.R8qYlc{-moz-border-radius:2px;border-radius:2px;background-color:rgba(97,97,97,0.902);position:absolute;left:0;width:100%;height:100%;opacity:0;transform:scale(0,0.5);transform-origin:inherit}.AZnilc{display:block;position:relative;font-size:10px;font-weight:500;padding:5px 8px 6px;opacity:0}.RM9ulf.qs41qe .R8qYlc{opacity:1;transform:scale(1,1)}.RM9ulf.catR2e .AZnilc{word-wrap:break-word}.RM9ulf.qs41qe .AZnilc{opacity:1}.RM9ulf.AXm5jc .AZnilc{font-size:14px;padding:8px 16px}.RM9ulf.u5lFJe{transition-property:-webkit-transform;transition-property:transform;transition-property:transform,-webkit-transform;transition-duration:200ms;transition-timing-function:cubic-bezier(0.24,1,0.32,1)}.RM9ulf.u5lFJe .R8qYlc{transition-property:opacity,-webkit-transform;transition-property:opacity,transform;transition-property:opacity,transform,-webkit-transform;transition-duration:50ms,200ms;transition-timing-function:linear,cubic-bezier(0.24,1,0.32,1)}.RM9ulf.u5lFJe .AZnilc{transition-property:opacity;transition-duration:150ms;transition-delay:50ms;transition-timing-function:cubic-bezier(0,0,0.6,1)}.RM9ulf.xCxor{transition-property:opacity;transition-duration:70ms;transition-delay:0ms;transition-timing-function:linear}sentinel{}</style><style id="vjrRq" nonce="">.ReaRCe{}</style><style nonce="" type="text/css" data-late-css="">.TYHMlb{display:block}.d3Fkdd.d3Fkdd.d3Fkdd{padding:0}.gKkZCe{align-items:center;border-bottom:0.0625rem solid #e0e0e0;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;padding:0.5rem 1rem}.yoswQd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.SNYuNc{box-flex:1;flex-grow:1;margin-left:1rem}.KeAbHb{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:0 1rem}.NyxV9b{justify-content:space-between;max-width:35rem;width:100%}.najF6d{margin-top:1rem;max-width:35rem}.zaxms{box-sizing:border-box;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;margin-top:1rem;padding:1.5rem}.Hc4hZd{margin-bottom:1rem}.iewtrc{max-width:100%;width:17.5rem}.U4xB8d{align-items:flex-start;box-sizing:border-box;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;margin:1rem;max-width:35rem;padding:0 1.5rem;width:100%}.U4xB8d ul{list-style:disc;margin-top:0.5rem;padding-left:1rem}.U4xB8d li{padding-bottom:1rem}.sH5Xkb{display:inline}sentinel{}</style><style nonce="" type="text/css" data-late-css="">.X5qqgf{max-width:35rem;overflow:visible;width:100%}.X5qqgf .wnIM7{overflow:initial}.HjNdme:not(:empty),.X5qqgf .yDGClf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-bottom:1rem}.VZ92zf{background-color:#d50000;color:#fff;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;font-size:0.8125rem;justify-content:space-between;line-height:1.25rem;margin:0.0625rem 0.0625rem;min-height:1.25rem;padding:0.5rem 1rem}.fyExH{background-color:#f5f5f5;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-top:1.5rem;overflow:hidden;padding:1rem}.asMx5b{margin:0}.W8M4Ad{margin-left:0.5rem}sentinel{}</style><style nonce="" type="text/css" data-late-css="">.RFWSze,.OkyLBb .oJeWuf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;overflow:hidden;justify-content:center}.OkyLBb .oJeWuf>.RFWSze,.RFWSze>.RFWSze{box-flex:1;flex-grow:1}.QngqV{margin:1rem 0}.OkyLBb .oJeWuf{margin-top:-1rem;padding:0;width:19.5rem}@media (min-height:HR_320_REM){.OkyLBb .oJeWuf{min-height:22.875rem}}.OkyLBb [role="separator"]{margin:0}.OkyLBb .aZsqhc{flex-shrink:0;padding:0.75rem 1.5rem}.hmmgFc,.Wsx9cf{margin:0.25rem 0;padding:1rem 1.5rem}.aZsqhc{flex-shrink:0;padding:1rem 1.5rem}.aZsqhc.RDPZE{opacity:.5}.s8kmpb{padding-left:1.5rem;padding-top:1rem}.GRzDxf{overflow:auto}.URRowe{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-right:2rem}sentinel{}</style><style nonce="" type="text/css" data-late-css="">.vgIUH{margin-bottom:1.25rem;text-align:center}.qDHZC{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:500}@media not all and (max-width:40rem){.FXCSf{min-width:25rem}}.picker-dialog.XKSfm-Sx9Kwc{-moz-box-shadow:rgba(0,0,0,.2) 0 0.25rem 1rem;box-shadow:rgba(0,0,0,.2) 0 0.25rem 1rem;background:#fff;-moz-box-shadow:0 0.25rem 1rem rgba(0,0,0,.12),0 0 0.25rem rgba(0,0,0,.12);box-shadow:0 0.25rem 1rem rgba(0,0,0,.12),0 0 0.25rem rgba(0,0,0,.12);padding:0;position:absolute;z-index:1194}.fFW7wc.XKSfm-Sx9Kwc{padding:0}.fFW7wc.XKSfm-Sx9Kwc-bN97Pc{border:0;height:23.125rem;margin:0;padding:0;position:relative;width:44.0625rem}.fFW7wc.XKSfm-Sx9Kwc-xJ5Hnf{background:#000;left:0;position:absolute;top:0;z-index:1193}.fFW7wc.XKSfm-Sx9Kwc-r4nke,.fFW7wc.XKSfm-Sx9Kwc-c6xFrd{display:none}.fFW7wc-OEVmcd{border:0;height:100%;overflow:hidden;width:100%}sentinel{}</style><link type="image/png" rel="icon" href="https://ssl.gstatic.com/classroom/favicon_black.png"><link type="image/png" rel="icon" href="https://ssl.gstatic.com/classroom/favicon_black.png"><link type="image/png" rel="icon" href="https://ssl.gstatic.com/classroom/favicon_black.png"><link type="image/png" rel="icon" href="https://ssl.gstatic.com/classroom/favicon_black.png"><style nonce="" type="text/css" data-late-css="">.yYWAMb{background:var(--dt-background,#fff);color:var(--dt-on-background,rgb(60,64,67))}.XV0XSd{--dt-display-1-font:400 4rem/4.75rem "Google Sans Display";--dt-display-1-spacing:0;--dt-display-large-font:400 3.5rem/4rem "Google Sans Display";--dt-display-large-spacing:0;--dt-display-medium-font:400 2.75rem/3.25rem "Google Sans Display";--dt-display-medium-spacing:0;--dt-display-small-font:400 2.25rem/2.75rem "Google Sans";--dt-display-small-spacing:0;--dt-headline-large-font:400 2rem/2.5rem "Google Sans";--dt-headline-large-spacing:0;--dt-headline-medium-font:400 1.75rem/2.25rem "Google Sans";--dt-headline-medium-spacing:0;--dt-headline-small-font:400 1.5rem/2rem "Google Sans";--dt-headline-small-spacing:0;--dt-title-large-font:400 1.375rem/1.75rem "Google Sans";--dt-title-large-spacing:0;--dt-headline-6-font:400 1.125rem/1.5rem "Google Sans";--dt-headline-6-spacing:0;--dt-title-medium-font:500 1rem/1.5rem "Google Sans";--dt-title-medium-spacing:0.00625em;--dt-title-small-font:500 0.875rem/1.25rem "Google Sans";--dt-title-small-spacing:0.0178571429em;--dt-subtitle-1-font:500 1rem/1.5rem "Roboto";--dt-subtitle-1-spacing:0.0125em;--dt-label-large-font:500 0.875rem/1.25rem "Roboto";--dt-label-large-spacing:0.0178571429em;--dt-label-medium-font:500 0.75rem/1rem "Roboto";--dt-label-medium-spacing:0.0208333333em;--dt-label-small-font:500 0.6875rem/1rem "Roboto";--dt-label-small-spacing:0.0727272727em;--dt-label-small-transform:uppercase;--dt-body-large-font:400 1rem/1.5rem "Roboto";--dt-body-large-spacing:0.00625em;--dt-body-medium-font:400 0.875rem/1.25rem "Roboto";--dt-body-medium-spacing:0.0142857143em;--dt-body-small-font:400 0.75rem/1rem "Roboto";--dt-body-small-spacing:0.025em;--dt-corner-banner:0.25rem;--dt-corner-button:0.25rem;--dt-corner-card:0.375rem;--dt-corner-card-thumbnail:0;--dt-corner-chip:6.25rem;--dt-corner-chip-avatar:6.25rem;--dt-corner-chip-suggestive:0.5rem;--dt-corner-dialog:0.5rem;--dt-corner-dialog-anchored:0.5rem;--dt-corner-fab:6.25rem;--dt-corner-fab-large:6.25rem;--dt-corner-field:0.375rem;--dt-corner-field-filled:0.375rem 0.375rem 0 0;--dt-corner-field-search:0.5rem;--dt-corner-icon-button:6.25rem;--dt-corner-landmark:0;--dt-corner-menu:0.25rem;--dt-corner-mole:0.25rem;--dt-corner-nav-drawer:0 1.5rem 1.5rem 0;--dt-corner-region:0.5rem;--dt-corner-tile:0.375rem}.vhoiae,.X9XeLb,.cWKK1c,.aJfoSc,.TOb6Ze{--dt-display-1-font:400 3.5625rem/4rem "Google Sans";--dt-display-1-spacing:0;--dt-display-large-font:400 3.5625rem/4rem "Google Sans";--dt-display-large-spacing:0;--dt-display-medium-font:400 2.8125rem/3.25rem "Google Sans";--dt-display-medium-spacing:0;--dt-display-small-font:400 2.25rem/2.75rem "Google Sans";--dt-display-small-spacing:0;--dt-headline-large-font:400 2rem/2.5rem "Google Sans";--dt-headline-large-spacing:0;--dt-headline-medium-font:400 1.75rem/2.25rem "Google Sans";--dt-headline-medium-spacing:0;--dt-headline-small-font:400 1.5rem/2rem "Google Sans";--dt-headline-small-spacing:0;--dt-title-large-font:400 1.375rem/1.75rem "Google Sans";--dt-title-large-spacing:0;--dt-headline-6-font:400 1.375rem/1.75rem "Google Sans";--dt-headline-6-spacing:0;--dt-title-medium-font:500 1rem/1.5rem "Google Sans Text";--dt-title-medium-spacing:0;--dt-title-small-font:500 0.875rem/1.25rem "Google Sans Text";--dt-title-small-spacing:0;--dt-subtitle-1-font:500 1rem/1.5rem "Google Sans Text";--dt-subtitle-1-spacing:0;--dt-label-large-font:500 0.875rem/1.25rem "Google Sans Text";--dt-label-large-spacing:0;--dt-label-medium-font:500 0.75rem/1rem "Google Sans Text";--dt-label-medium-spacing:0;--dt-label-small-font:500 0.6875rem/1rem "Google Sans Text";--dt-label-small-spacing:0.0090909091em;--dt-label-small-transform:none;--dt-body-large-font:400 1rem/1.5rem "Google Sans Text";--dt-body-large-spacing:0;--dt-body-medium-font:400 0.875rem/1.25rem "Google Sans Text";--dt-body-medium-spacing:0;--dt-body-small-font:400 0.75rem/1rem "Google Sans Text";--dt-body-small-spacing:0.0083333333em;--dt-corner-banner:0.5rem;--dt-corner-button:6.25rem;--dt-corner-card:0.75rem;--dt-corner-card-thumbnail:0.25rem;--dt-corner-chip:0.5rem;--dt-corner-chip-avatar:6.25rem;--dt-corner-chip-suggestive:0.5rem;--dt-corner-dialog:0.5rem;--dt-corner-dialog-anchored:0.5rem;--dt-corner-fab:1rem;--dt-corner-fab-large:1.75rem;--dt-corner-field:0.25rem;--dt-corner-field-filled:0.25rem 0.25rem 0 0;--dt-corner-field-search:0.25rem;--dt-corner-icon-button:6.25rem;--dt-corner-landmark:1rem;--dt-corner-menu:0.25rem;--dt-corner-mole:1rem;--dt-corner-nav-drawer:6.25rem;--dt-corner-region:0.75rem;--dt-corner-tile:1rem;scrollbar-width:8px;scrollbar-color:var(--dt-outline-variant,rgb(218,220,224)) transparent}.vhoiae .tk3N6e-suEOdc,.X9XeLb .tk3N6e-suEOdc,.cWKK1c .tk3N6e-suEOdc,.aJfoSc .tk3N6e-suEOdc,.TOb6Ze .tk3N6e-suEOdc{font:var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-small-spacing,.025em);background:var(--dt-inverse-surface,rgb(32,33,36));border-radius:.25rem;border:solid 1px transparent;-moz-box-sizing:border-box;box-sizing:border-box;color:var(--dt-inverse-on-surface,rgb(218,220,224));margin:0;max-width:100vw;min-height:1.375rem;min-width:3.5rem;padding:.25rem .5rem;text-align:center;z-index:6000}.vhoiae .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd),.X9XeLb .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd),.cWKK1c .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd),.aJfoSc .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd),.TOb6Ze .tk3N6e-suEOdc:not(.tk3N6e-suEOdc-ZYIfFd){opacity:1;transform:scale(1);transition:opacity 45ms linear,transform .15s _tooltip_transform_easing}.vhoiae .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd,.X9XeLb .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd,.cWKK1c .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd,.aJfoSc .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd,.TOb6Ze .tk3N6e-suEOdc.tk3N6e-suEOdc-ZYIfFd{opacity:0;transform:scale(.9);width:0}.vhoiae .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo,.X9XeLb .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo,.cWKK1c .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo,.aJfoSc .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo,.TOb6Ze .tk3N6e-suEOdc .tk3N6e-suEOdc-hFsbo{display:none}.vhoiae .XKSfm-Sx9Kwc,.X9XeLb .XKSfm-Sx9Kwc,.cWKK1c .XKSfm-Sx9Kwc,.aJfoSc .XKSfm-Sx9Kwc,.TOb6Ze .XKSfm-Sx9Kwc{background-color:var(--dt-surface,#fff);border-radius:var(--dt-corner-dialog,.5rem);color:var(--dt-on-surface,rgb(60,64,67))}.vhoiae .XKSfm-Sx9Kwc-bN97Pc,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,.0142857143em);background-color:var(--dt-surface,#fff)}.vhoiae .XKSfm-Sx9Kwc-r4nke,.X9XeLb .XKSfm-Sx9Kwc-r4nke,.cWKK1c .XKSfm-Sx9Kwc-r4nke,.aJfoSc .XKSfm-Sx9Kwc-r4nke,.TOb6Ze .XKSfm-Sx9Kwc-r4nke{background-color:var(--dt-surface,#fff)}.vhoiae .XKSfm-Sx9Kwc-r4nke-TvD9Pc,.X9XeLb .XKSfm-Sx9Kwc-r4nke-TvD9Pc,.cWKK1c .XKSfm-Sx9Kwc-r4nke-TvD9Pc,.aJfoSc .XKSfm-Sx9Kwc-r4nke-TvD9Pc,.TOb6Ze .XKSfm-Sx9Kwc-r4nke-TvD9Pc{color:var(--dt-on-surface,rgb(60,64,67))}.vhoiae .XKSfm-Sx9Kwc-r4nke-fmcmS,.X9XeLb .XKSfm-Sx9Kwc-r4nke-fmcmS,.cWKK1c .XKSfm-Sx9Kwc-r4nke-fmcmS,.aJfoSc .XKSfm-Sx9Kwc-r4nke-fmcmS,.TOb6Ze .XKSfm-Sx9Kwc-r4nke-fmcmS{font:var(--dt-headline-small-font,400 1.5rem/2rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-headline-small-spacing,0)}.vhoiae .XKSfm-Sx9Kwc-dI4VCc,.X9XeLb .XKSfm-Sx9Kwc-dI4VCc,.cWKK1c .XKSfm-Sx9Kwc-dI4VCc,.aJfoSc .XKSfm-Sx9Kwc-dI4VCc,.TOb6Ze .XKSfm-Sx9Kwc-dI4VCc{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,.0142857143em);background-color:var(--dt-surface,#fff);border-color:var(--dt-outline,rgb(128,134,139));border-radius:var(--dt-corner-field,.375rem);-moz-box-sizing:border-box;box-sizing:border-box;color:var(--dt-on-surface,rgb(60,64,67));height:2.625rem}.vhoiae .XKSfm-Sx9Kwc-dI4VCc:focus,.X9XeLb .XKSfm-Sx9Kwc-dI4VCc:focus,.cWKK1c .XKSfm-Sx9Kwc-dI4VCc:focus,.aJfoSc .XKSfm-Sx9Kwc-dI4VCc:focus,.TOb6Ze .XKSfm-Sx9Kwc-dI4VCc:focus{border-color:var(--dt-primary,rgb(26,115,232));border-width:.125rem;box-shadow:none}.vhoiae .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc,.X9XeLb .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc,.cWKK1c .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc,.aJfoSc .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc,.TOb6Ze .euCgFf-CJXtmf-Sx9Kwc .XKSfm-Sx9Kwc-bN97Pc{background:none}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe{font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,.0178571429em);overflow:visible;border-radius:var(--dt-corner-button,.25rem);color:var(--dt-primary,rgb(26,115,232));text-transform:capitalize}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button::after,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe::after{transition:color 15ms linear,background 15ms linear,opacity 15ms linear}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:active,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:hover,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:active,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:hover,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:active,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:hover,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:active,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:hover,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:active,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:hover,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:active,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:hover,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:active,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:hover,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:active,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:hover,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:active,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:hover,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:active,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:hover,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover{box-shadow:none}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before{background-color:currentcolor}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::before{border-radius:var(--dt-corner-button,.25rem);opacity:.12}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:hover::before{border-radius:var(--dt-corner-button,.25rem);opacity:.08}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button:focus::after,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button:focus::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button:focus::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button:focus::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button:focus::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button:focus::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button:focus::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button:focus::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe:focus::after{bottom:0;border-radius:.375rem;content:"";display:block;height:100%;left:0;outline:solid 2px var(--dt-primary,rgb(26,115,232));outline-offset:3px;position:absolute;width:100%}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc{overflow:visible;background-color:var(--dt-primary,rgb(26,115,232));color:var(--dt-on-primary,#fff)}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc::after{transition:color 15ms linear,background 15ms linear,opacity 15ms linear}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover{box-shadow:none}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before{background-color:currentcolor}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::before{border-radius:var(--dt-corner-button,.25rem);opacity:.12}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:hover::before{border-radius:var(--dt-corner-button,.25rem);opacity:.08}.vhoiae .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc button.VIpgJd-ldDVFe-JIbuQc:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd button.VIpgJd-ldDVFe-JIbuQc:focus::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.VIpgJd-ldDVFe-JIbuQc:focus::after{bottom:0;border-radius:.375rem;content:"";display:block;height:100%;left:0;outline:solid 2px var(--dt-primary,rgb(26,115,232));outline-offset:3px;position:absolute;width:100%}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe{padding-top:.3125rem}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc{background-color:var(--dt-surface,#fff);background-image:none;border:.0625rem solid var(--dt-outline,rgb(128,134,139));box-shadow:none;-moz-box-sizing:border-box;box-sizing:border-box;color:var(--dt-primary,rgb(26,115,232))}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:active,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:focus,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:hover{border:.0625rem solid var(--dt-outline,rgb(128,134,139));box-shadow:none}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me){overflow:visible}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me),.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me)::after{transition:color 15ms linear,background 15ms linear,opacity 15ms linear}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover{box-shadow:none}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before{background-color:currentcolor}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::before{border-radius:var(--dt-corner-button,.25rem);opacity:.12}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):hover::before{border-radius:var(--dt-corner-button,.25rem);opacity:.08}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc:not(.tk3N6e-LgbsSe-OWB6Me):focus::after{bottom:0;border-radius:.375rem;content:"";display:block;height:100%;left:0;outline:solid 2px var(--dt-primary,rgb(26,115,232));outline-offset:3px;position:absolute;width:100%}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me{color:var(--dt-on-background,rgb(60,64,67));opacity:.38}.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.vhoiae .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.vhoiae .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.X9XeLb .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.X9XeLb .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.cWKK1c .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.cWKK1c .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.aJfoSc .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.aJfoSc .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-bN97Pc .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:active::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:focus::before,.TOb6Ze .XKSfm-Sx9Kwc-c6xFrd .tk3N6e-LgbsSe.tk3N6e-LgbsSe-haDnnc.tk3N6e-LgbsSe-OWB6Me:hover::before{background-color:inherit}.vhoiae ::-webkit-scrollbar,.X9XeLb ::-webkit-scrollbar,.cWKK1c ::-webkit-scrollbar,.aJfoSc ::-webkit-scrollbar,.TOb6Ze ::-webkit-scrollbar{height:8px;width:8px}.vhoiae ::-webkit-scrollbar-corner,.X9XeLb ::-webkit-scrollbar-corner,.cWKK1c ::-webkit-scrollbar-corner,.aJfoSc ::-webkit-scrollbar-corner,.TOb6Ze ::-webkit-scrollbar-corner{background:transparent}.vhoiae ::-webkit-scrollbar-thumb,.X9XeLb ::-webkit-scrollbar-thumb,.cWKK1c ::-webkit-scrollbar-thumb,.aJfoSc ::-webkit-scrollbar-thumb,.TOb6Ze ::-webkit-scrollbar-thumb{background-clip:padding-box;background-color:var(--dt-outline-variant,rgb(218,220,224));border-radius:100px;border:none;height:8px;padding:100px 0 0;width:8px}.vhoiae ::-webkit-scrollbar-thumb:hover,.X9XeLb ::-webkit-scrollbar-thumb:hover,.cWKK1c ::-webkit-scrollbar-thumb:hover,.aJfoSc ::-webkit-scrollbar-thumb:hover,.TOb6Ze ::-webkit-scrollbar-thumb:hover{background-color:var(--dt-outline,rgb(128,134,139))}.vhoiae ::-webkit-scrollbar-thumb:active,.X9XeLb ::-webkit-scrollbar-thumb:active,.cWKK1c ::-webkit-scrollbar-thumb:active,.aJfoSc ::-webkit-scrollbar-thumb:active,.TOb6Ze ::-webkit-scrollbar-thumb:active{background-color:var(--dt-outline,rgb(128,134,139))}.vhoiae ::-webkit-scrollbar-track,.X9XeLb ::-webkit-scrollbar-track,.cWKK1c ::-webkit-scrollbar-track,.aJfoSc ::-webkit-scrollbar-track,.TOb6Ze ::-webkit-scrollbar-track{background-color:transparent;border:none;box-shadow:none;height:8px;width:8px}.vhoiae ::-webkit-scrollbar-track:hover,.X9XeLb ::-webkit-scrollbar-track:hover,.cWKK1c ::-webkit-scrollbar-track:hover,.aJfoSc ::-webkit-scrollbar-track:hover,.TOb6Ze ::-webkit-scrollbar-track:hover{border:none;box-shadow:none}@media (forced-colors:active){.vhoiae ::-webkit-scrollbar-thumb,.vhoiae ::-webkit-scrollbar-thumb:hover,.vhoiae ::-webkit-scrollbar-thumb:active,.X9XeLb ::-webkit-scrollbar-thumb,.X9XeLb ::-webkit-scrollbar-thumb:hover,.X9XeLb ::-webkit-scrollbar-thumb:active,.cWKK1c ::-webkit-scrollbar-thumb,.cWKK1c ::-webkit-scrollbar-thumb:hover,.cWKK1c ::-webkit-scrollbar-thumb:active,.aJfoSc ::-webkit-scrollbar-thumb,.aJfoSc ::-webkit-scrollbar-thumb:hover,.aJfoSc ::-webkit-scrollbar-thumb:active,.TOb6Ze ::-webkit-scrollbar-thumb,.TOb6Ze ::-webkit-scrollbar-thumb:hover,.TOb6Ze ::-webkit-scrollbar-thumb:active{background-color:CanvasText}}.XV0XSd.KkxPLb{--dt-background:#fff;--dt-on-background:rgb(60,64,67);--dt-on-background-secondary:rgb(95,99,104);--dt-outline:rgb(128,134,139);--dt-outline-variant:rgb(218,220,224);--dt-on-disabled:rgba(60,64,67,0.38);--dt-disabled:rgba(60,64,67,0.12);--dt-inverse-on-surface:rgb(218,220,224);--dt-inverse-surface:rgb(32,33,36);--dt-on-surface-variant:rgb(95,99,104);--dt-on-surface-secondary:rgb(95,99,104);--dt-on-surface:rgb(60,64,67);--dt-surface-tint:rgb(241,243,244);--dt-surface-variant:rgb(241,243,244);--dt-surface1:#fff;--dt-surface1-shadow:0 1px 2px 0 rgba(60,64,67,0.3),0 1px 3px 1px rgba(60,64,67,0.15);--dt-surface2:#fff;--dt-surface2-shadow:0 1px 2px 0 rgba(60,64,67,0.3),0 2px 6px 2px rgba(60,64,67,0.15);--dt-surface3:#fff;--dt-surface3-shadow:0 1px 3px 0 rgba(60,64,67,0.3),0 4px 8px 3px rgba(60,64,67,0.15);--dt-surface4:#fff;--dt-surface4-shadow:0 2px 3px 0 rgba(60,64,67,0.3),0 6px 10px 4px rgba(60,64,67,0.15);--dt-surface5:#fff;--dt-surface5-shadow:0 4px 4px 0 rgba(60,64,67,0.3),0 8px 12px 6px rgba(60,64,67,0.15);--dt-surface:#fff;--dt-scrim:rgba(32,33,36,0.6);--dt-scrim-2x:rgb(32,33,36);--dt-on-primary-container:rgb(60,64,67);--dt-on-primary:#fff;--dt-primary-action-state-layer:rgb(25,103,210);--dt-primary-action-stateful:rgb(24,90,188);--dt-primary-action:rgb(25,103,210);--dt-primary-container-icon:rgb(25,103,210);--dt-primary-container-link:rgb(25,103,210);--dt-primary-container:rgb(232,240,254);--dt-primary-icon:#fff;--dt-primary-link:#fff;--dt-primary-outline:rgb(24,90,188);--dt-primary:rgb(26,115,232);--dt-on-secondary-container:rgb(60,64,67);--dt-on-secondary:#fff;--dt-secondary-action-state-layer:rgb(60,64,67);--dt-secondary-action-stateful:rgb(32,33,36);--dt-secondary-action:rgb(60,64,67);--dt-secondary-container-icon:rgb(60,64,67);--dt-secondary-container-link:rgb(25,103,210);--dt-secondary-container:rgb(241,243,244);--dt-secondary-icon:#fff;--dt-secondary-link:#fff;--dt-secondary-outline:rgb(60,64,67);--dt-secondary:rgb(60,64,67);--dt-on-tertiary-container:rgb(60,64,67);--dt-on-tertiary:#fff;--dt-tertiary-action-state-layer:rgb(19,115,51);--dt-tertiary-action-stateful:rgb(13,101,45);--dt-tertiary-action:rgb(19,115,51);--dt-tertiary-container-icon:rgb(19,115,51);--dt-tertiary-container-link:rgb(19,115,51);--dt-tertiary-container:rgb(230,244,234);--dt-tertiary-icon:#fff;--dt-tertiary-link:#fff;--dt-tertiary-outline:rgb(19,115,51);--dt-tertiary:rgb(24,128,56);--dt-on-neutral-container:rgb(60,64,67);--dt-on-neutral:#fff;--dt-neutral-action-state-layer:rgb(60,64,67);--dt-neutral-action-stateful:rgb(32,33,36);--dt-neutral-action:rgb(60,64,67);--dt-neutral-container-icon:rgb(60,64,67);--dt-neutral-container-link:rgb(25,103,210);--dt-neutral-container:rgb(241,243,244);--dt-neutral-icon:#fff;--dt-neutral-link:#fff;--dt-neutral-outline:rgb(60,64,67);--dt-neutral:rgb(60,64,67);--dt-error-action-state-layer:rgb(197,34,31);--dt-error-action-stateful:rgb(179,20,18);--dt-error-action:rgb(197,34,31);--dt-error-container-icon:rgb(197,34,31);--dt-error-container-link:rgb(197,34,31);--dt-error-container:rgb(252,232,230);--dt-error-icon:#fff;--dt-error-link:#fff;--dt-error-outline:rgb(179,20,18);--dt-error:rgb(217,48,37);--dt-on-error-container:rgb(60,64,67);--dt-on-error:#fff;--dt-on-warning-container:rgb(60,64,67);--dt-on-warning:rgb(32,33,36);--dt-warning-action-state-layer:rgb(234,134,0);--dt-warning-action-stateful:rgb(32,33,36);--dt-warning-action:rgb(60,64,67);--dt-warning-container-icon:rgb(60,64,67);--dt-warning-container-link:rgb(60,64,67);--dt-warning-container:rgb(254,247,224);--dt-warning-icon:rgb(60,64,67);--dt-warning-link:rgb(60,64,67);--dt-warning-outline:rgb(234,134,0);--dt-warning:rgb(249,171,0)}.XV0XSd.LgGVmb{--dt-background:rgb(32,33,36);--dt-on-background:rgb(232,234,237);--dt-on-background-secondary:rgb(154,160,166);--dt-outline:rgb(95,99,104);--dt-outline-variant:rgb(189,193,198);--dt-on-disabled:rgba(232,234,237,0.38);--dt-disabled:rgba(232,234,237,0.12);--dt-inverse-on-surface:rgb(60,64,67);--dt-inverse-surface:rgb(241,243,244);--dt-on-surface-secondary:rgb(154,160,166);--dt-on-surface-variant:rgb(154,160,166);--dt-on-surface:rgb(232,234,237);--dt-surface-tint:rgb(60,64,67);--dt-surface-variant:rgb(60,64,67);--dt-surface1:rgb(32,33,36);--dt-surface1-shadow:0 1px 2px 0 rgba(0,0,0,0.3),0 1px 3px 1px rgba(0,0,0,0.15);--dt-surface2:rgb(32,33,36);--dt-surface2-shadow:0 1px 2px 0 rgba(0,0,0,0.3),0 2px 6px 2px rgba(0,0,0,0.15);--dt-surface3:#36373a;--dt-surface3-shadow:0 1px 3px 0 rgba(0,0,0,0.3),0 4px 8px 3px rgba(0,0,0,0.15);--dt-surface4:rgb(32,33,36);--dt-surface4-shadow:0 2px 3px 0 rgba(0,0,0,0.3),0 6px 10px 4px rgba(0,0,0,0.15);--dt-surface5:rgb(32,33,36);--dt-surface5-shadow:0 4px 4px 0 rgba(0,0,0,0.3),0 8px 12px 6px rgba(0,0,0,0.15);--dt-surface:rgb(32,33,36);--dt-scrim:rgba(32,33,36,0.87);--dt-scrim-2x:rgb(241,243,244);--dt-on-primary-container:rgb(210,227,252);--dt-on-primary:rgb(32,33,36);--dt-primary-action-state-layer:rgb(138,180,248);--dt-primary-action-stateful:rgb(174,203,250);--dt-primary-action:rgb(138,180,248);--dt-primary-container-icon:rgb(210,227,252);--dt-primary-container-link:rgb(210,227,252);--dt-primary-container:#394457;--dt-primary-icon:rgb(32,33,36);--dt-primary-link:rgb(32,33,36);--dt-primary-outline:rgb(138,180,248);--dt-primary:rgb(138,180,248);--dt-on-secondary-container:rgb(241,243,244);--dt-on-secondary:rgb(218,220,224);--dt-secondary-action-state-layer:rgb(218,220,224);--dt-secondary-action-stateful:rgb(232,234,237);--dt-secondary-action:rgb(218,220,224);--dt-secondary-container-icon:rgb(241,243,244);--dt-secondary-container-link:rgb(241,243,244);--dt-secondary-container:#4d4e51;--dt-secondary-icon:rgb(218,220,224);--dt-secondary-link:rgb(218,220,224);--dt-secondary-outline:rgb(218,220,224);--dt-secondary:rgb(32,33,36);--dt-on-tertiary-container:rgb(206,234,214);--dt-on-tertiary:rgb(32,33,36);--dt-tertiary-action-state-layer:rgb(129,201,149);--dt-tertiary-action-stateful:rgb(168,218,181);--dt-tertiary-action:rgb(129,201,149);--dt-tertiary-container-icon:rgb(206,234,214);--dt-tertiary-container-link:rgb(206,234,214);--dt-tertiary-container:#37493f;--dt-tertiary-icon:rgb(32,33,36);--dt-tertiary-link:rgb(32,33,36);--dt-tertiary-outline:rgb(129,201,149);--dt-tertiary:rgb(129,201,149);--dt-on-neutral-container:rgb(232,234,237);--dt-on-neutral:rgb(32,33,36);--dt-neutral-action-state-layer:rgb(232,234,237);--dt-neutral-action-stateful:#fff;--dt-neutral-action:rgb(232,234,237);--dt-neutral-container-icon:rgb(232,234,237);--dt-neutral-container-link:rgb(174,203,250);--dt-neutral-container:rgb(60,64,67);--dt-neutral-icon:rgb(32,33,36);--dt-neutral-link:rgb(32,33,36);--dt-neutral-outline:rgb(232,234,237);--dt-neutral:rgb(232,234,237);--dt-error-action-state-layer:rgb(242,139,130);--dt-error-action-stateful:rgb(246,174,169);--dt-error-action:rgb(242,139,130);--dt-error-container-icon:rgb(250,210,207);--dt-error-container-link:rgb(250,210,207);--dt-error-container:#523a3b;--dt-error-icon:rgb(32,33,36);--dt-error-link:rgb(32,33,36);--dt-error-outline:rgb(242,139,130);--dt-error:rgb(242,139,130);--dt-on-error-container:rgb(250,210,207);--dt-on-error:rgb(32,33,36);--dt-on-warning-container:rgb(254,239,195);--dt-on-warning:rgb(32,33,36);--dt-warning-action-state-layer:rgb(253,214,99);--dt-warning-action-stateful:rgb(253,226,147);--dt-warning-action:rgb(253,214,99);--dt-warning-container-icon:rgb(254,239,195);--dt-warning-container-link:rgb(254,239,195);--dt-warning-container:#554c33;--dt-warning-icon:rgb(32,33,36);--dt-warning-link:rgb(32,33,36);--dt-warning-outline:rgb(253,214,99);--dt-warning:rgb(253,214,99)}.vhoiae.KkxPLb{--dt-on-background:#1F1F1F;--dt-on-background-secondary:#5E5E5E;--dt-background:#FFF;--dt-on-surface:#1F1F1F;--dt-inverse-surface:#303030;--dt-on-surface-secondary:#5E5E5E;--dt-on-surface-variant:#444746;--dt-surface-variant:#E3E3E3;--dt-inverse-on-surface:#F2F2F2;--dt-surface:#FFF;--dt-surface-tint:#6991d6;--dt-surface1:#f7f9fc;--dt-surface1-shadow:0px 3px 1px -2px rgba(0,0,0,0.2),0px 2px 2px 0px rgba(0,0,0,0.14),0px 1px 5px 0px rgba(0,0,0,0.12);--dt-surface2:#f2f6fc;--dt-surface2-shadow:0px 2px 4px -1px rgba(0,0,0,0.2),0px 4px 5px 0px rgba(0,0,0,0.14),0px 1px 10px 0px rgba(0,0,0,0.12);--dt-surface3:#edf2fc;--dt-surface3-shadow:0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12);--dt-surface4:#e8effb;--dt-surface4-shadow:0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12);--dt-surface5:#e2ecfb;--dt-surface5-shadow:0px 8px 10px -6px rgba(0,0,0,0.2),0px 16px 24px 2px rgba(0,0,0,0.14),0px 6px 30px 5px rgba(0,0,0,0.12);--dt-scrim:rgba(0,0,0,0.32);--dt-scrim-2x:rgba(0,0,0,0.64);--dt-on-primary-container:#041E49;--dt-primary-container-icon:#041E49;--dt-primary-container-link:#041E49;--dt-primary:#0B57D0;--dt-primary-action:#0B57D0;--dt-primary-action-stateful:#0B57D0;--dt-primary-outline:#0B57D0;--dt-primary-action-state-layer:#0B57D0;--dt-primary-container:#D3E3FD;--dt-on-primary:#FFF;--dt-primary-icon:#FFF;--dt-primary-link:#FFF;--dt-on-secondary-container:#001D35;--dt-secondary-container-icon:#001D35;--dt-secondary-container-link:#001D35;--dt-secondary:#00639B;--dt-secondary-action:#00639B;--dt-secondary-action-stateful:#00639B;--dt-secondary-outline:#00639B;--dt-secondary-action-state-layer:#00639B;--dt-secondary-container:#C2E7FF;--dt-on-secondary:#FFF;--dt-secondary-icon:#FFF;--dt-secondary-link:#FFF;--dt-on-tertiary-container:#072711;--dt-tertiary-container-icon:#072711;--dt-tertiary-container-link:#072711;--dt-tertiary:#146C2E;--dt-tertiary-action:#146C2E;--dt-tertiary-action-stateful:#146C2E;--dt-tertiary-outline:#146C2E;--dt-tertiary-action-state-layer:#146C2E;--dt-tertiary-container:#C4EED0;--dt-on-tertiary:#FFF;--dt-tertiary-icon:#FFF;--dt-tertiary-link:#FFF;--dt-on-neutral-container:#1F1F1F;--dt-neutral-container-icon:#1F1F1F;--dt-neutral-container-link:#1F1F1F;--dt-neutral:#474747;--dt-neutral-action:#1F1F1F;--dt-neutral-action-stateful:#1F1F1F;--dt-neutral-outline:#1F1F1F;--dt-neutral-action-state-layer:#1F1F1F;--dt-neutral-container:#E3E3E3;--dt-on-neutral:#FFF;--dt-neutral-icon:#FFF;--dt-neutral-link:#FFF;--dt-on-warning-container:#421F00;--dt-warning-container-icon:#421F00;--dt-warning-container-link:#421F00;--dt-warning:#F09D00;--dt-warning-action:#421F00;--dt-warning-action-stateful:#421F00;--dt-warning-outline:#421F00;--dt-warning-action-state-layer:#421F00;--dt-warning-container:#FFDF99;--dt-on-warning:#1F1F1F;--dt-warning-icon:#1F1F1F;--dt-warning-link:#1F1F1F;--dt-on-error-container:#410E0B;--dt-error-container-icon:#410E0B;--dt-error-container-link:#410E0B;--dt-error:#B3261E;--dt-error-action:#B3261E;--dt-error-action-stateful:#B3261E;--dt-error-outline:#B3261E;--dt-error-action-state-layer:#B3261E;--dt-error-container:#F9DEDC;--dt-on-error:#FFF;--dt-error-icon:#FFF;--dt-error-link:#FFF;--dt-disabled:rgba(31,31,31,0.12);--dt-on-disabled:rgba(31,31,31,0.38);--dt-outline:#747775;--dt-outline-variant:#C7C7C7}.vhoiae.LgGVmb{--dt-on-background:#E3E3E3;--dt-on-background-secondary:#ABABAB;--dt-background:#1F1F1F;--dt-on-surface:#E3E3E3;--dt-inverse-surface:#E3E3E3;--dt-on-surface-secondary:#ABABAB;--dt-on-surface-variant:#C4C7C5;--dt-surface-variant:#444746;--dt-inverse-on-surface:#303030;--dt-surface:#1F1F1F;--dt-surface-tint:#d1e1ff;--dt-surface1:#292a2d;--dt-surface1-shadow:0px 3px 1px -2px rgba(0,0,0,0.2),0px 2px 2px 0px rgba(0,0,0,0.14),0px 1px 5px 0px rgba(0,0,0,0.12);--dt-surface2:#2d2f33;--dt-surface2-shadow:0px 2px 4px -1px rgba(0,0,0,0.2),0px 4px 5px 0px rgba(0,0,0,0.14),0px 1px 10px 0px rgba(0,0,0,0.12);--dt-surface3:#31343a;--dt-surface3-shadow:0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12);--dt-surface4:#32363c;--dt-surface4-shadow:0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12);--dt-surface5:#353940;--dt-surface5-shadow:0px 8px 10px -6px rgba(0,0,0,0.2),0px 16px 24px 2px rgba(0,0,0,0.14),0px 6px 30px 5px rgba(0,0,0,0.12);--dt-scrim:rgba(0,0,0,0.32);--dt-scrim-2x:rgba(0,0,0,0.64);--dt-on-primary-container:#D3E3FD;--dt-primary-container-icon:#D3E3FD;--dt-primary-container-link:#D3E3FD;--dt-primary:#A8C7FA;--dt-primary-action:#A8C7FA;--dt-primary-action-stateful:#A8C7FA;--dt-primary-outline:#A8C7FA;--dt-primary-action-state-layer:#1B6EF3;--dt-primary-container:#0842A0;--dt-on-primary:#062E6F;--dt-primary-icon:#062E6F;--dt-primary-link:#062E6F;--dt-on-secondary-container:#C2E7FF;--dt-secondary-container-icon:#C2E7FF;--dt-secondary-container-link:#C2E7FF;--dt-secondary:#7FCFFF;--dt-secondary-action:#7FCFFF;--dt-secondary-action-stateful:#7FCFFF;--dt-secondary-outline:#7FCFFF;--dt-secondary-action-state-layer:#047DB7;--dt-secondary-container:#004A77;--dt-on-secondary:#035;--dt-secondary-icon:#035;--dt-secondary-link:#035;--dt-on-tertiary-container:#C4EED0;--dt-tertiary-container-icon:#C4EED0;--dt-tertiary-container-link:#C4EED0;--dt-tertiary:#6DD58C;--dt-tertiary-action:#6DD58C;--dt-tertiary-action-stateful:#6DD58C;--dt-tertiary-outline:#6DD58C;--dt-tertiary-action-state-layer:#198639;--dt-tertiary-container:#0F5223;--dt-on-tertiary:#0A3818;--dt-tertiary-icon:#0A3818;--dt-tertiary-link:#0A3818;--dt-on-neutral-container:#E3E3E3;--dt-neutral-container-icon:#E3E3E3;--dt-neutral-container-link:#E3E3E3;--dt-neutral:#ABABAB;--dt-neutral-action:#ABABAB;--dt-neutral-action-stateful:#ABABAB;--dt-neutral-outline:#ABABAB;--dt-neutral-action-state-layer:#ABABAB;--dt-neutral-container:#474747;--dt-on-neutral:#1F1F1F;--dt-neutral-icon:#ABABAB;--dt-neutral-link:#ABABAB;--dt-on-warning-container:#FFF0D1;--dt-warning-container-icon:#FFF0D1;--dt-warning-container-link:#FFF0D1;--dt-warning:#FFBB29;--dt-warning-action:#FFBB29;--dt-warning-action-stateful:#FFBB29;--dt-warning-outline:#FFF0D1;--dt-warning-action-state-layer:#FFBB29;--dt-warning-container:#562D00;--dt-on-warning:#1F1F1F;--dt-warning-icon:#421F00;--dt-warning-link:#421F00;--dt-on-error-container:#F9DEDC;--dt-error-container-icon:#F9DEDC;--dt-error-container-link:#F9DEDC;--dt-error:#F2B8B5;--dt-error-action:#F2B8B5;--dt-error-action-stateful:#F2B8B5;--dt-error-outline:#F2B8B5;--dt-error-action-state-layer:#DC362E;--dt-error-container:#8C1D18;--dt-on-error:#601410;--dt-error-icon:#601410;--dt-error-link:#601410;--dt-disabled:rgba(227,227,227,0.12);--dt-on-disabled:rgba(227,227,227,0.38);--dt-outline:#8E918F;--dt-outline-variant:#444746}.XV0XSd .yYWAMb.bvmRsc,.XV0XSd .dif24c.bvmRsc{--dt-background:rgb(32,33,36);--dt-on-background:rgb(232,234,237);--dt-on-background-secondary:rgb(154,160,166);--dt-outline:rgb(95,99,104);--dt-outline-variant:rgb(189,193,198);--dt-on-disabled:rgba(232,234,237,0.38);--dt-disabled:rgba(232,234,237,0.12);--dt-inverse-on-surface:rgb(60,64,67);--dt-inverse-surface:rgb(241,243,244);--dt-on-surface-secondary:rgb(154,160,166);--dt-on-surface-variant:rgb(154,160,166);--dt-on-surface:rgb(232,234,237);--dt-surface-tint:rgb(60,64,67);--dt-surface-variant:rgb(60,64,67);--dt-surface1:rgb(32,33,36);--dt-surface1-shadow:0 1px 2px 0 rgba(0,0,0,0.3),0 1px 3px 1px rgba(0,0,0,0.15);--dt-surface2:rgb(32,33,36);--dt-surface2-shadow:0 1px 2px 0 rgba(0,0,0,0.3),0 2px 6px 2px rgba(0,0,0,0.15);--dt-surface3:#36373a;--dt-surface3-shadow:0 1px 3px 0 rgba(0,0,0,0.3),0 4px 8px 3px rgba(0,0,0,0.15);--dt-surface4:rgb(32,33,36);--dt-surface4-shadow:0 2px 3px 0 rgba(0,0,0,0.3),0 6px 10px 4px rgba(0,0,0,0.15);--dt-surface5:rgb(32,33,36);--dt-surface5-shadow:0 4px 4px 0 rgba(0,0,0,0.3),0 8px 12px 6px rgba(0,0,0,0.15);--dt-surface:rgb(32,33,36);--dt-scrim:rgba(32,33,36,0.87);--dt-scrim-2x:rgb(241,243,244);--dt-on-primary-container:rgb(210,227,252);--dt-on-primary:rgb(32,33,36);--dt-primary-action-state-layer:rgb(138,180,248);--dt-primary-action-stateful:rgb(174,203,250);--dt-primary-action:rgb(138,180,248);--dt-primary-container-icon:rgb(210,227,252);--dt-primary-container-link:rgb(210,227,252);--dt-primary-container:#394457;--dt-primary-icon:rgb(32,33,36);--dt-primary-link:rgb(32,33,36);--dt-primary-outline:rgb(138,180,248);--dt-primary:rgb(138,180,248);--dt-on-secondary-container:rgb(241,243,244);--dt-on-secondary:rgb(218,220,224);--dt-secondary-action-state-layer:rgb(218,220,224);--dt-secondary-action-stateful:rgb(232,234,237);--dt-secondary-action:rgb(218,220,224);--dt-secondary-container-icon:rgb(241,243,244);--dt-secondary-container-link:rgb(241,243,244);--dt-secondary-container:#4d4e51;--dt-secondary-icon:rgb(218,220,224);--dt-secondary-link:rgb(218,220,224);--dt-secondary-outline:rgb(218,220,224);--dt-secondary:rgb(32,33,36);--dt-on-tertiary-container:rgb(206,234,214);--dt-on-tertiary:rgb(32,33,36);--dt-tertiary-action-state-layer:rgb(129,201,149);--dt-tertiary-action-stateful:rgb(168,218,181);--dt-tertiary-action:rgb(129,201,149);--dt-tertiary-container-icon:rgb(206,234,214);--dt-tertiary-container-link:rgb(206,234,214);--dt-tertiary-container:#37493f;--dt-tertiary-icon:rgb(32,33,36);--dt-tertiary-link:rgb(32,33,36);--dt-tertiary-outline:rgb(129,201,149);--dt-tertiary:rgb(129,201,149);--dt-on-neutral-container:rgb(232,234,237);--dt-on-neutral:rgb(32,33,36);--dt-neutral-action-state-layer:rgb(232,234,237);--dt-neutral-action-stateful:#fff;--dt-neutral-action:rgb(232,234,237);--dt-neutral-container-icon:rgb(232,234,237);--dt-neutral-container-link:rgb(174,203,250);--dt-neutral-container:rgb(60,64,67);--dt-neutral-icon:rgb(32,33,36);--dt-neutral-link:rgb(32,33,36);--dt-neutral-outline:rgb(232,234,237);--dt-neutral:rgb(232,234,237);--dt-error-action-state-layer:rgb(242,139,130);--dt-error-action-stateful:rgb(246,174,169);--dt-error-action:rgb(242,139,130);--dt-error-container-icon:rgb(250,210,207);--dt-error-container-link:rgb(250,210,207);--dt-error-container:#523a3b;--dt-error-icon:rgb(32,33,36);--dt-error-link:rgb(32,33,36);--dt-error-outline:rgb(242,139,130);--dt-error:rgb(242,139,130);--dt-on-error-container:rgb(250,210,207);--dt-on-error:rgb(32,33,36);--dt-on-warning-container:rgb(254,239,195);--dt-on-warning:rgb(32,33,36);--dt-warning-action-state-layer:rgb(253,214,99);--dt-warning-action-stateful:rgb(253,226,147);--dt-warning-action:rgb(253,214,99);--dt-warning-container-icon:rgb(254,239,195);--dt-warning-container-link:rgb(254,239,195);--dt-warning-container:#554c33;--dt-warning-icon:rgb(32,33,36);--dt-warning-link:rgb(32,33,36);--dt-warning-outline:rgb(253,214,99);--dt-warning:rgb(253,214,99)}.vhoiae .yYWAMb.bvmRsc,.vhoiae .dif24c.bvmRsc,.X9XeLb .yYWAMb.bvmRsc,.X9XeLb .dif24c.bvmRsc,.cWKK1c .yYWAMb.bvmRsc,.cWKK1c .dif24c.bvmRsc,.aJfoSc .yYWAMb.bvmRsc,.aJfoSc .dif24c.bvmRsc,.TOb6Ze .yYWAMb.bvmRsc,.TOb6Ze .dif24c.bvmRsc{--dt-on-background:#E3E3E3;--dt-on-background-secondary:#ABABAB;--dt-background:#1F1F1F;--dt-on-surface:#E3E3E3;--dt-inverse-surface:#E3E3E3;--dt-on-surface-secondary:#ABABAB;--dt-on-surface-variant:#C4C7C5;--dt-surface-variant:#444746;--dt-inverse-on-surface:#303030;--dt-surface:#1F1F1F;--dt-surface-tint:#d1e1ff;--dt-surface1:#292a2d;--dt-surface1-shadow:0px 3px 1px -2px rgba(0,0,0,0.2),0px 2px 2px 0px rgba(0,0,0,0.14),0px 1px 5px 0px rgba(0,0,0,0.12);--dt-surface2:#2d2f33;--dt-surface2-shadow:0px 2px 4px -1px rgba(0,0,0,0.2),0px 4px 5px 0px rgba(0,0,0,0.14),0px 1px 10px 0px rgba(0,0,0,0.12);--dt-surface3:#31343a;--dt-surface3-shadow:0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12);--dt-surface4:#32363c;--dt-surface4-shadow:0px 5px 5px -3px rgba(0,0,0,0.2),0px 8px 10px 1px rgba(0,0,0,0.14),0px 3px 14px 2px rgba(0,0,0,0.12);--dt-surface5:#353940;--dt-surface5-shadow:0px 8px 10px -6px rgba(0,0,0,0.2),0px 16px 24px 2px rgba(0,0,0,0.14),0px 6px 30px 5px rgba(0,0,0,0.12);--dt-scrim:rgba(0,0,0,0.32);--dt-scrim-2x:rgba(0,0,0,0.64);--dt-on-primary-container:#D3E3FD;--dt-primary-container-icon:#D3E3FD;--dt-primary-container-link:#D3E3FD;--dt-primary:#A8C7FA;--dt-primary-action:#A8C7FA;--dt-primary-action-stateful:#A8C7FA;--dt-primary-outline:#A8C7FA;--dt-primary-action-state-layer:#1B6EF3;--dt-primary-container:#0842A0;--dt-on-primary:#062E6F;--dt-primary-icon:#062E6F;--dt-primary-link:#062E6F;--dt-on-secondary-container:#C2E7FF;--dt-secondary-container-icon:#C2E7FF;--dt-secondary-container-link:#C2E7FF;--dt-secondary:#7FCFFF;--dt-secondary-action:#7FCFFF;--dt-secondary-action-stateful:#7FCFFF;--dt-secondary-outline:#7FCFFF;--dt-secondary-action-state-layer:#047DB7;--dt-secondary-container:#004A77;--dt-on-secondary:#035;--dt-secondary-icon:#035;--dt-secondary-link:#035;--dt-on-tertiary-container:#C4EED0;--dt-tertiary-container-icon:#C4EED0;--dt-tertiary-container-link:#C4EED0;--dt-tertiary:#6DD58C;--dt-tertiary-action:#6DD58C;--dt-tertiary-action-stateful:#6DD58C;--dt-tertiary-outline:#6DD58C;--dt-tertiary-action-state-layer:#198639;--dt-tertiary-container:#0F5223;--dt-on-tertiary:#0A3818;--dt-tertiary-icon:#0A3818;--dt-tertiary-link:#0A3818;--dt-on-neutral-container:#E3E3E3;--dt-neutral-container-icon:#E3E3E3;--dt-neutral-container-link:#E3E3E3;--dt-neutral:#ABABAB;--dt-neutral-action:#ABABAB;--dt-neutral-action-stateful:#ABABAB;--dt-neutral-outline:#ABABAB;--dt-neutral-action-state-layer:#ABABAB;--dt-neutral-container:#474747;--dt-on-neutral:#1F1F1F;--dt-neutral-icon:#ABABAB;--dt-neutral-link:#ABABAB;--dt-on-warning-container:#FFF0D1;--dt-warning-container-icon:#FFF0D1;--dt-warning-container-link:#FFF0D1;--dt-warning:#FFBB29;--dt-warning-action:#FFBB29;--dt-warning-action-stateful:#FFBB29;--dt-warning-outline:#FFF0D1;--dt-warning-action-state-layer:#FFBB29;--dt-warning-container:#562D00;--dt-on-warning:#1F1F1F;--dt-warning-icon:#421F00;--dt-warning-link:#421F00;--dt-on-error-container:#F9DEDC;--dt-error-container-icon:#F9DEDC;--dt-error-container-link:#F9DEDC;--dt-error:#F2B8B5;--dt-error-action:#F2B8B5;--dt-error-action-stateful:#F2B8B5;--dt-error-outline:#F2B8B5;--dt-error-action-state-layer:#DC362E;--dt-error-container:#8C1D18;--dt-on-error:#601410;--dt-error-icon:#601410;--dt-error-link:#601410;--dt-disabled:rgba(227,227,227,0.12);--dt-on-disabled:rgba(227,227,227,0.38);--dt-outline:#8E918F;--dt-outline-variant:#444746}.Q6yead{fill:currentcolor;overflow:hidden}.mig17c{overflow:visible}[dir=rtl] .Q6yead.wSyMnf{transform:scaleX(-1)}@media (forced-colors:active){.Q6yead.QJZfhe.QJZfhe{fill:CanvasText}}.A5Gtre{font:inherit;font-size:100%;font-weight:inherit;text-decoration:none}.A5Gtre:hover,.A5Gtre:active,.A5Gtre:focus{text-decoration:underline}.cS0c5e{clip-path:inset(50%);clip:rect(1px,1px,1px,1px);height:1px;margin:-1px;opacity:0;overflow:hidden;padding:0;position:absolute;width:1px}.tk3N6e-VCkuzd{-moz-box-shadow:0 1px 3px rgba(0,0,0,.2);box-shadow:0 1px 3px rgba(0,0,0,.2);background-color:#fff;border:1px solid;border-color:#bbb #bbb #a8a8a8;padding:16px;position:absolute;z-index:1201!important}.tk3N6e-VCkuzd-hFsbo{position:absolute}.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc,.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG{display:block;height:0;position:absolute;width:0}.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-jQ8oHc{border:9px solid}.tk3N6e-VCkuzd-hFsbo .tk3N6e-VCkuzd-ez0xG{border:8px solid}.tk3N6e-VCkuzd-Ya1KTb{bottom:0}.tk3N6e-VCkuzd-d6mlqf{top:-9px}.tk3N6e-VCkuzd-y6n2Me{left:-9px}.tk3N6e-VCkuzd-cX0Lwc{right:0}.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc{left:-9px}.tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc{border-color:#bbb transparent;left:-9px}.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc{border-color:#a8a8a8 transparent}.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-ez0xG,.tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-ez0xG{border-color:#fff transparent;left:-8px}.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-jQ8oHc,.tk3N6e-VCkuzd-Ya1KTb .tk3N6e-VCkuzd-ez0xG{border-bottom-width:0}.tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-jQ8oHc{border-top-width:0}.tk3N6e-VCkuzd-d6mlqf .tk3N6e-VCkuzd-ez0xG{border-top-width:0;top:1px}.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-jQ8oHc,.tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-jQ8oHc{border-color:transparent #bbb;top:-9px}.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-ez0xG,.tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-ez0xG{border-color:transparent #fff;top:-8px}.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-jQ8oHc{border-left-width:0}.tk3N6e-VCkuzd-y6n2Me .tk3N6e-VCkuzd-ez0xG{border-left-width:0;left:1px}.tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-jQ8oHc,.tk3N6e-VCkuzd-cX0Lwc .tk3N6e-VCkuzd-ez0xG{border-right-width:0}.tk3N6e-suEOdc{-moz-border-radius:0;border-radius:0;-moz-box-shadow:none;box-shadow:none;-moz-transition:visibility 0,opacity 0.13s ease-in;transition:visibility 0,opacity 0.13s ease-in;background-color:#2a2a2a;border:1px solid #fff;color:#fff;cursor:default;display:block;font-size:11px;font-weight:bold;margin-left:-1px;opacity:1;padding:7px 9px;position:absolute;visibility:visible;white-space:pre-wrap;word-break:break-all;word-break:break-word}.tk3N6e-suEOdc-ZYIfFd{-moz-transition:visibility 0.13s,opacity 0.13s ease-out,left 0 linear 0.13s,top 0 linear 0.13s;transition:visibility 0.13s,opacity 0.13s ease-out,left 0 linear 0.13s,top 0 linear 0.13s;opacity:0;left:20px!important;top:20px!important;visibility:hidden}.tk3N6e-suEOdc-wZVHld{display:none}.tk3N6e-suEOdc-hFsbo{pointer-events:none;position:absolute}.tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc,.tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG{content:"";display:block;height:0;position:absolute;width:0}.tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-jQ8oHc{border:6px solid}.tk3N6e-suEOdc-hFsbo .tk3N6e-suEOdc-ez0xG{border:5px solid}.tk3N6e-suEOdc-Ya1KTb{bottom:0}.tk3N6e-suEOdc-d6mlqf{top:-6px}.tk3N6e-suEOdc-y6n2Me{left:-6px}.tk3N6e-suEOdc-cX0Lwc{right:0}.tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc,.tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc{border-color:#fff transparent;left:-6px}.tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG,.tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG{border-color:#2a2a2a transparent;left:-5px}.tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc,.tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG{border-bottom-width:0}.tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc{border-top-width:0}.tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG{border-top-width:0;top:1px}.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc,.tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc{border-color:transparent #fff;top:-6px}.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG,.tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG{border-color:transparent #2a2a2a;top:-5px}.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc{border-left-width:0}.tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG{border-left-width:0;left:1px}.tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc,.tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG{border-right-width:0}.cAHxfe{font:var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-small-spacing,.025em);background:var(--dt-inverse-surface,rgb(32,33,36));border-radius:.25rem;border:solid 1px transparent;-moz-box-sizing:border-box;box-sizing:border-box;color:var(--dt-inverse-on-surface,rgb(218,220,224));margin:0;max-width:100vw;min-height:1.375rem;min-width:3.5rem;padding:.25rem .5rem;text-align:center;z-index:6000}.cAHxfe:not(.tk3N6e-suEOdc-ZYIfFd){opacity:1;transform:scale(1);transition:opacity 45ms linear,transform .15s _tooltip_transform_easing}.cAHxfe.tk3N6e-suEOdc-ZYIfFd{opacity:0;transform:scale(.9);width:0}.cAHxfe .tk3N6e-suEOdc-hFsbo{display:none}.pDtC4e{display:inline-block}@keyframes shimmer{0%{background-position:100% 50%}to{background-position:0 50%}}@keyframes fadeInAnimation{0%{opacity:0}to{opacity:1}}.ja0jmf{align-content:center;animation-fill-mode:forwards;animation-iteration-count:1;animation:fadeInAnimation ease 200ms;background-color:var(--dt-surface,#fff);display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;height:100%;position:absolute;top:0;width:100%;z-index:3000}.F6wkof{animation:shimmer 2.2s ease infinite;background:0 0/300% 300% linear-gradient(-61deg,var(--dt-inverse-on-surface,#dadce0) 40%,var(--dt-surface-variant,#f1f3f4) 50%,var(--dt-inverse-on-surface,#dadce0) 60%);background-color:var(--dt-inverse-on-surface,#dadce0)}@media (forced-colors:active){.F6wkof{border:1px solid var(--dt-outline,#80868b)}}.HrDxdd{-moz-border-radius:1rem;border-radius:1rem;height:1rem;margin-left:1rem;margin-top:.5rem}.HrDxdd:nth-child(odd){margin-top:1.5rem}.ISv2N{background-color:transparent;border:none;color:inherit;cursor:pointer;fill:currentColor;margin-right:1rem;margin-top:.125rem;outline:none;padding:.75rem;text-decoration:none}.EebkFb{align-items:center;border-bottom:1px solid var(--dt-outline,#80868b);display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:space-between;margin-bottom:1rem;margin-top:.3125rem;padding-bottom:.375rem;width:100%}.gAm2E{font:var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-title-medium-spacing,0.00625em);color:var(--dt-on-background,#3c4043);margin-left:20px}.NFRm8d{align-items:center;animation-fill-mode:forwards;animation-iteration-count:1;animation:fadeInAnimation ease 200ms;background-color:var(--dt-surface,#fff);display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;height:100%;width:100%;z-index:3000}.C4MDDc{font:var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-small-spacing,0.025em);color:var(--dt-on-surface,#3c4043);margin-top:5.125rem}@media (forced-colors:active){.RCmsv{background-color:ButtonFace!important}.RCmsv,.RCmsv::before{border-color:ButtonText!important}.RCmsv:disabled,.RCmsv.RDPZE,.RCmsv:disabled::before,.RCmsv.RDPZE::before{border-color:GrayText!important;opacity:1!important}.RCmsv.u3bW4e,.RCmsv:focus,.RCmsv:hover,.hp3b6d.u3bW4e,.hp3b6d:focus,.hp3b6d:hover{background-color:Highlight!important}.RCmsv.u3bW4e,.RCmsv:focus,.RCmsv:hover,.hp3b6d.u3bW4e,.hp3b6d:focus,.hp3b6d:hover,.RCmsv.u3bW4e::before,.RCmsv:focus::before,.RCmsv:hover::before,.hp3b6d.u3bW4e::before,.hp3b6d:focus::before,.hp3b6d:hover::before{border-color:HighlightText!important;outline-color:HighlightText!important}.jbArdc,.jbArdc [viewBox]{color:ButtonText!important;fill:currentcolor!important;forced-color-adjust:none}.jbArdc:disabled,.jbArdc.RDPZE,.jbArdc:disabled [viewBox],.jbArdc.RDPZE [viewBox]{color:GrayText!important;opacity:1!important}.jbArdc.u3bW4e,.jbArdc:focus,.jbArdc:hover,.jbArdc.u3bW4e [viewBox],.jbArdc:focus [viewBox],.jbArdc:hover [viewBox]{color:HighlightText!important}.Yz4sEb{background-color:Field!important;border-color:FieldText!important}.Yz4sEb:disabled,.Yz4sEb.RDPZE{border-color:GrayText!important}.GyDQo{color:FieldText!important;fill:currentcolor!important;forced-color-adjust:none}.GyDQo:disabled,.GyDQo.RDPZE{color:GrayText!important;opacity:1!important}.GyDQo::-webkit-input-placeholder{color:GrayText!important;opacity:1!important}.GyDQo::-moz-placeholder{color:GrayText!important;opacity:1!important}.GyDQo:-ms-input-placeholder{color:GrayText!important;opacity:1!important}.GyDQo::-ms-input-placeholder{color:GrayText!important;opacity:1!important}.GyDQo::placeholder{color:GrayText!important;opacity:1!important}.cNqOse{background-color:Canvas!important}.cNqOse.kUXOd{border-color:CanvasText!important;border-style:solid!important;border-width:1px!important}.X0gZEc{color:CanvasText!important;fill:currentcolor!important;forced-color-adjust:none}.ObwPwb{background-color:Highlight!important}.rkFgee{color:HighlightText!important;fill:currentcolor!important;forced-color-adjust:none}.uevTLb{color:LinkText!important;fill:currentcolor!important;forced-color-adjust:none}.uevTLb:active,.uevTLb.qs41qe{color:ActiveText!important}.uevTLb:visited,.uevTLb.gxDgLe{color:VisitedText!important}}.I1PgQd{-moz-box-sizing:border-box;box-sizing:border-box;padding:.5rem 1rem;width:20rem}.ousvBd{-moz-box-align:center;align-items:center;display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-right:-.5rem}.Zcp8g.vKmmhc{color:var(--dt-on-surface,#3c4043);font-size:1.25rem;line-height:1.25rem;margin-right:.3rem}.nCnYNd{font:var(--dt-title-small-font,500 .875rem/1.25rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-title-small-spacing,0.0178571429em);color:var(--dt-on-surface,#3c4043);-moz-box-flex:1;-moz-box-flex:1;flex:1}.EafEFe{font:var(--dt-title-large-font,400 1.375rem/1.75rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-title-large-spacing,0);margin-bottom:.75rem}.RQM9Gf{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em);color:var(--dt-on-surface,#3c4043)}.EIsVy{display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-pack:end;justify-content:flex-end;margin:0 -.25rem}.BjbK3c{border-width:0;box-shadow:0px 1px 2px 0px rgba(60,64,67,.30),0px 2px 6px 2px rgba(60,64,67,.15);background:var(--dt-surface2,#fff);-moz-border-radius:.5rem;border-radius:.5rem;position:relative}.BjbK3c::before{border:solid 1px transparent;-moz-border-radius:inherit;border-radius:inherit;bottom:0;content:"";left:0;position:absolute;right:0;top:0}.kaZy8e,.cDqddf,.FfqPSe,.kAgEFc{fill:var(--dt-background,#fff);position:absolute}.kaZy8e,.FfqPSe{height:1.0625rem;left:50%;margin-left:-0.9375rem;width:1.875rem}.kaZy8e{top:-1.0625rem}.FfqPSe{bottom:-1.0625rem}.cDqddf,.kAgEFc{height:1.875rem;margin-top:-0.9375rem;top:50%;width:1.0625rem}.cDqddf{right:-1.0625rem}.kAgEFc{left:-1.0625rem}.ob9sLd{font:var(--dt-body-small-font,400 .75rem/1rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-small-spacing,.025em);border-radius:.25rem;-moz-box-sizing:border-box;box-sizing:border-box;display:inline-block;font-weight:500;height:1.25rem;line-height:1.25rem;overflow:hidden;padding:0 .5rem;position:relative;text-overflow:ellipsis;white-space:nowrap}.ob9sLd::before{border:solid 1px transparent;border-radius:inherit;bottom:0;content:"";left:0;position:absolute;right:0;top:0}@media (forced-colors:active){.ob9sLd::before{border-color:CanvasText}}.Chn84b-haAclf{left:0;top:0;background-color:transparent;border:none;height:100%;width:100%;overflow:hidden;padding:0;position:absolute;z-index:2500}.Chn84b-haAclf.xTMeO{display:none}.Chn84b-L5Fo6c-haAclf{height:100%;width:100%;background:transparent;padding:0;position:absolute;z-index:1}.ge6pde .Chn84b-L5Fo6c-haAclf{opacity:0}.Chn84b-o1DAbe-aZ2wEe-Lb81de{-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%);left:50%;position:absolute;top:50%;z-index:1}.Chn84b-o1DAbe-ge6pde-haAclf-Lb81de{position:absolute;left:0;right:0;top:0;bottom:0;overflow:hidden;border:none;padding:0;display:-webkit-box;display:-webkit-flex;display:-moz-box;display:-ms-flexbox;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;-moz-box-align:center;align-items:center;-moz-box-pack:center;justify-content:center;background-color:rgba(32,33,36,.6);visibility:hidden;z-index:2}.ge6pde .Chn84b-o1DAbe-ge6pde-haAclf-Lb81de{visibility:visible}.Chn84b-o1DAbe-ge6pde-Sx9Kwc-Lb81de{width:616px;height:516px;max-width:616px;max-height:516px;min-width:512px;min-height:272px;-moz-border-radius:8px;border-radius:8px;background-color:white;padding:0;margin:20px;overflow:hidden;position:relative}.Chn84b-o1DAbe-ge6pde-fmcmS-Lb81de{color:rgba(32,33,36,.87);font-size:22px;left:24px;position:absolute;top:26px}.Chn84b-o1DAbe-ge6pde-TvD9Pc-LgbsSe{background:url(https://fonts.gstatic.com/s/i/short-term/release/googlesymbols/close/default/24px.svg);border:0;cursor:pointer;height:24px;opacity:.87;position:absolute;right:24px;top:22px;width:24px}.Chn84b-o1DAbe-ge6pde-TvD9Pc-suEOdc{visibility:hidden;-moz-border-radius:2px;border-radius:2px;border:0;background-color:#202124;color:#fff;position:absolute;z-index:1;right:24px;top:48px;opacity:1;overflow-x:hidden;padding:5px 8px 6px;text-align:center;font-size:12px}.Chn84b-o1DAbe-ge6pde-TvD9Pc:hover .Chn84b-o1DAbe-ge6pde-TvD9Pc-suEOdc{visibility:visible}.oErxNe-pSzOP{width:36px;height:36px;overflow:hidden;-moz-animation:mspin-rotate 1568.63ms infinite linear}.oErxNe-pSzOP .oErxNe-WkJb5{-moz-animation:mspin-revrot 5332ms infinite steps(4)}.oErxNe-pSzOP .oErxNe-aZ2wEe{background-image:url("//ssl.gstatic.com/docs/picker/images/loading_spinner.svg");background-size:100%;width:11664px;height:36px;-moz-animation:mspin-medium-film 5332ms infinite steps(324)}@keyframes mspin-medium-film{0%{transform:translateX(0)}to{transform:translateX(-11664px)}}@keyframes mspin-rotate{0%{transform:rotate(0deg)}to{transform:rotate(360deg)}}@keyframes mspin-revrot{0%{transform:rotate(0deg)}to{transform:rotate(-360deg)}}@keyframes mspin-medium-film{0%{transform:translateX(0)}to{transform:translateX(-11664px)}}.ndfHFb-aZ2wEe{height:44px;overflow:hidden;position:relative}.ndfHFb-vyDMJf-aZ2wEe{height:28px;left:50%;margin-left:-14px;position:absolute;top:8px;width:28px}.ndfHFb-vyDMJf-aZ2wEe.auswjd{animation:container-rotate 1568ms linear infinite}@keyframes container-rotate{to{transform:rotate(360deg)}}.aZ2wEe-pbTTYe{position:absolute;width:100%;height:100%;opacity:0}.aZ2wEe-v3pZbf{border-color:#4285f4}.aZ2wEe-oq6NAc{border-color:#db4437}.aZ2wEe-gS7Ybc{border-color:#f4b400}.aZ2wEe-nllRtd{border-color:#0f9d58}.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-v3pZbf{animation:fill-unfill-rotate 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both,blue-fade-in-out 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both}.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-oq6NAc{animation:fill-unfill-rotate 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both,red-fade-in-out 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both}.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-gS7Ybc{animation:fill-unfill-rotate 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both,yellow-fade-in-out 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both}.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-pbTTYe.aZ2wEe-nllRtd{animation:fill-unfill-rotate 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both,green-fade-in-out 5332ms cubic-bezier(0.4,0.0,0.2,1) infinite both}@keyframes fill-unfill-rotate{12.5%{transform:rotate(135deg)}25%{transform:rotate(270deg)}37.5%{transform:rotate(405deg)}50%{transform:rotate(540deg)}62.5%{transform:rotate(675deg)}75%{transform:rotate(810deg)}87.5%{transform:rotate(945deg)}to{transform:rotate(1080deg)}}@keyframes blue-fade-in-out{0%{opacity:1}25%{opacity:1}26%{opacity:0}89%{opacity:0}90%{opacity:1}to{opacity:1}}@keyframes red-fade-in-out{0%{opacity:0}15%{opacity:0}25%{opacity:1}50%{opacity:1}51%{opacity:0}}@keyframes yellow-fade-in-out{0%{opacity:0}40%{opacity:0}50%{opacity:1}75%{opacity:1}76%{opacity:0}}@keyframes green-fade-in-out{0%{opacity:0}65%{opacity:0}75%{opacity:1}90%{opacity:1}to{opacity:0}}.aZ2wEe-pehrl-TpMipd{position:absolute;box-sizing:border-box;top:0;left:45%;width:10%;height:100%;overflow:hidden;border-color:inherit}.aZ2wEe-pehrl-TpMipd .aZ2wEe-LkdAo{width:1000%;left:-450%}.aZ2wEe-LkdAo-e9ayKc{display:inline-block;position:relative;width:50%;height:100%;overflow:hidden;border-color:inherit}.aZ2wEe-LkdAo-e9ayKc .aZ2wEe-LkdAo{width:200%}.aZ2wEe-LkdAo{box-sizing:border-box;height:100%;border-width:3px;border-style:solid;border-color:inherit;border-bottom-color:transparent!important;-moz-border-radius:50%;border-radius:50%;animation:none}.aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo{border-right-color:transparent!important;transform:rotate(129deg)}.aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo{left:-100%;border-left-color:transparent!important;transform:rotate(-129deg)}.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-LK5yu .aZ2wEe-LkdAo{animation:left-spin 1333ms cubic-bezier(0.4,0.0,0.2,1) infinite both}.ndfHFb-vyDMJf-aZ2wEe.auswjd .aZ2wEe-LkdAo-e9ayKc.aZ2wEe-qwU8Me .aZ2wEe-LkdAo{animation:right-spin 1333ms cubic-bezier(0.4,0.0,0.2,1) infinite both}@keyframes left-spin{0%{transform:rotate(130deg)}50%{transform:rotate(-5deg)}to{transform:rotate(130deg)}}@keyframes right-spin{0%{transform:rotate(-130deg)}50%{transform:rotate(5deg)}to{transform:rotate(-130deg)}}.aZ2wEe-hj4D6d{position:absolute;top:0;bottom:0;right:0;left:0}.wvGCSb-VkLyEc-Sx9Kwc{font-size:14px;white-space:normal;width:472px}.wvGCSb-VkLyEc-Sx9Kwc .wvGCSb-VkLyEc-Sx9Kwc-VdSJob{width:424px}.wvGCSb-VkLyEc-Sx9Kwc .HB1eCd-HzV7m-LgbsSe-bN97Pc{font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif}.wvGCSb{color:black;font-family:Arial,sans-serif,sans;font-family:var(--docs-material-font-family,Arial,sans-serif,sans);font-size:13px;white-space:normal}.wvGCSb.HB1eCd-UMrnmb{font-size:14px}.wvGCSb .tk3N6e-LgbsSe{font-family:Arial,sans-serif,sans;font-family:var(--docs-material-header-font-family,Arial,sans-serif,sans);font-weight:700;font-weight:var(--docs-material-font-weight-bold,700)}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe{margin:0 8px 0 0;min-width:24px;vertical-align:middle}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe-ZmdkE{box-shadow:none;background-color:rgba(0,0,0,.06);background-image:none;cursor:pointer;border-color:transparent!important;border-radius:2px;border-width:1px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe-auswjd{box-shadow:none;background-color:rgba(0,0,0,.12);background-image:none;cursor:pointer;border-color:transparent!important;border-radius:2px;border-width:1px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e{border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:white;border:1px solid #dadce0!important;color:#1a73e8;height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-OWB6Me{border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:white;border:1px solid #f1f3f4!important;color:#3c4043;opacity:.38;height:24px;padding:3px 12px 5px}@media (forced-colors:active){.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-XpnDCe{outline:1px solid Highlight;outline-offset:-4px}}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe{border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#e9f1fe;border:1px solid #c1d8fb!important;height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-ZmdkE{border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#f8fbff;border:1px solid #cce0fc!important;height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE{border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#e1ecfe;border:1px solid #bbd4fb!important;height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-n2to0e.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd{border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#e1ecfe;border:1px solid transparent!important;box-shadow:0 2px 6px 2px rgba(60,64,67,.15);height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc{background-image:none;border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#1a73e8;color:#fff;height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-OWB6Me{background-image:none;border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#1a73e8;color:#fff;background:#f8f9fa;color:#202124;opacity:.62;height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe{background-image:none;border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#1a73e8;color:#fff;background:#5094ed;box-shadow:0 1px 3px 1px rgba(66,133,244,.15);height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-ZmdkE{background-image:none;border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#1a73e8;color:#fff;background:#2b7de9;box-shadow:0 1px 3px 1px rgba(66,133,244,.15);height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-ZmdkE{background-image:none;border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#1a73e8;color:#fff;background:#63a0ef;box-shadow:0 1px 3px 1px rgba(66,133,244,.15);height:24px;padding:3px 12px 5px}.wvGCSb.HB1eCd-UMrnmb .tk3N6e-LgbsSe.tk3N6e-LgbsSe-JIbuQc.tk3N6e-LgbsSe-XpnDCe.tk3N6e-LgbsSe-auswjd{background-image:none;border:1px solid transparent!important;border-radius:4px;box-shadow:none;box-sizing:border-box;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-weight:500;font-size:14px;height:36px;letter-spacing:.25px;line-height:16px;padding:9px 24px 11px 24px;background:#1a73e8;color:#fff;background:#63a0ef;box-shadow:0 2px 6px 2px rgba(66,133,244,.15);height:24px;padding:3px 12px 5px}.wvGCSb .XKSfm-Sx9Kwc-c6xFrd{font-family:Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-family:var(--docs-material-header-font-family,Roboto,RobotoDraft,Helvetica,Arial,sans-serif);font-weight:500}.wvGCSb .XKSfm-Sx9Kwc-r4nke{font-size:16px}.HB1eCd-UMrnmb .wvGCSb .XKSfm-Sx9Kwc-r4nke{font-size:22px}.wvGCSb .XKSfm-Sx9Kwc-r4nke-fmcmS{font-family:Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-family:var(--docs-material-header-font-family,Roboto,RobotoDraft,Helvetica,Arial,sans-serif);font-weight:normal}.HB1eCd-UMrnmb .lI7fHe-XKSfm.XKSfm-Sx9Kwc{width:300px}.HB1eCd-UMrnmb .lI7fHe-XKSfm .XKSfm-Sx9Kwc-r4nke-fmcmS{display:block;width:220px;word-wrap:break-word}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc{background:#fff;border:1px solid transparent;border-radius:8px;box-shadow:0 4px 8px 3px rgba(60,64,67,.15);position:absolute;z-index:1003}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-xJ5Hnf{background-color:#000;left:0;position:absolute;top:0;z-index:998}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc:focus{outline:none}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke{border-bottom:none;padding:24px}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-fmcmS{color:#202124;font-family:"Google Sans",Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-size:22px;font-weight:400;line-height:28px}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-r4nke-TvD9Pc{height:24px;position:absolute;right:24px;top:26px;width:24px}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-bN97Pc{min-width:312px;padding:0 24px 24px;color:#3c4043;font-family:Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-size:13px;font-size:var(--docs-material-font-size-normal,13px)}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc-c6xFrd{display:flex;justify-content:flex-end;padding:24px}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc .HB1eCd-HzV7m-LgbsSe-edvN0e-ssJRIf.HB1eCd-HzV7m-LgbsSe{margin-left:12px;text-transform:none}.HB1eCd-HzV7m-UMrnmb-Sx9Kwc .HB1eCd-HzV7m-LgbsSe-aSvl1d-zTETae.HB1eCd-HzV7m-LgbsSe{text-transform:none}.ndfHFb-c4YZDc-Sx9Kwc{background:#fff;background-clip:padding-box;border:1px solid #acacac;border:1px solid rgba(0,0,0,.333);-moz-box-shadow:0 4px 16px rgba(0,0,0,.2);box-shadow:0 4px 16px rgba(0,0,0,.2);outline:0;padding:30px 42px;position:absolute;z-index:1195}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-Sx9Kwc{background:var(--dt-surface,#fff);padding:24px 24px;-moz-border-radius:8px;border-radius:8px}.ndfHFb-c4YZDc-Sx9Kwc-xJ5Hnf{background-color:#000;left:0;position:absolute;top:0;z-index:1194}.ndfHFb-c4YZDc-qbOKL-OEVmcd .VIpgJd-TUo6Hb-xJ5Hnf,.ndfHFb-c4YZDc-qbOKL-OEVmcd .XKSfm-Sx9Kwc-xJ5Hnf{background-color:#000}div.ndfHFb-c4YZDc-Sx9Kwc-xJ5Hnf{filter:alpha(opacity=75);opacity:.75}.ndfHFb-c4YZDc-Sx9Kwc-r4nke{background-color:#fff;color:#000;cursor:default;font-size:16px;line-height:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-r4nke{background-color:var(--dt-surface,#fff);color:var(--dt-on-surface,#3c4043);font:var(--dt-headline-small-font,400 1.5rem/2rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-headline-small-spacing,0)}.ndfHFb-c4YZDc-Sx9Kwc-r4nke-TvD9Pc{height:11px;filter:alpha(opacity=70);opacity:.7;padding:17px;position:absolute;right:0;top:0;width:11px}.ndfHFb-c4YZDc-Sx9Kwc-r4nke-TvD9Pc:after{content:"";background:url(//ssl.gstatic.com/ui/v1/dialog/close-x.png);position:absolute;height:11px;width:11px;right:17px}.ndfHFb-c4YZDc-Sx9Kwc-r4nke-TvD9Pc:hover{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-Sx9Kwc-bN97Pc{background-color:#fff;line-height:1.4em}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-bN97Pc{background-color:var(--dt-surface,#fff)}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button{-moz-border-radius:2px;border-radius:2px;background-color:#f5f5f5;background-image:-moz-linear-gradient(top,#f5f5f5,#f1f1f1);background-image:linear-gradient(top,#f5f5f5,#f1f1f1);border:1px solid #dcdcdc;border:1px solid rgba(0,0,0,.1);color:#444;cursor:default;font-size:11px;font-weight:bold;height:29px;line-height:27px;margin:0 16px 0 0;min-width:72px;outline:0;padding:0 8px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button{margin:0 0 0 24px;line-height:20px;-moz-border-radius:100px;border-radius:100px;background:var(--dt-surface,#fff);color:var(--dt-primary,#1a73e8);font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em);border:none}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:hover,.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:active{-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1);background-color:#f8f8f8;background-image:-moz-linear-gradient(top,#f8f8f8,#f1f1f1);background-image:linear-gradient(top,#f8f8f8,#f1f1f1);border:1px solid #c6c6c6;color:#333}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:hover{background:rgba(168,199,250,.08);color:var(--dt-primary,#1a73e8);border:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:focus,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:active{background:rgba(168,199,250,.12);color:var(--dt-primary,#1a73e8);border:none;outline:none;-moz-box-shadow:none;box-shadow:none}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:active{-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.1);box-shadow:inset 0 1px 2px rgba(0,0,0,.1)}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button:focus{border:1px solid #4d90fe}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd button[disabled]{-moz-box-shadow:none;box-shadow:none;background:#fff;background-image:none;border:1px solid #f3f3f3;border:1px solid rgba(0,0,0,.05);color:#b8b8b8}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc{background-color:#1a73e8;background-image:-moz-linear-gradient(top,#4d90fe,#4787ed);background-image:linear-gradient(top,#4d90fe,#4787ed);border:1px solid #3079ed;color:#fff}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc:hover{background-color:#357ae8;background-image:-moz-linear-gradient(top,#4d90fe,#357ae8);background-image:linear-gradient(top,#4d90fe,#357ae8);border:1px solid #2f5bb7;color:#fff}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc:active{background-color:#357ae8;background-image:-moz-linear-gradient(top,#4d90fe,#357ae8);background-image:linear-gradient(top,#4d90fe,#357ae8);border:1px solid #2f5bb7;color:#fff;-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.3);box-shadow:inset 0 1px 2px rgba(0,0,0,.3)}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc:focus{-moz-box-shadow:inset 0 0 0 1px #fff;box-shadow:inset 0 0 0 1px #fff;border:1px solid #fff;border:rgba(0,0,0,0) solid 1px;outline:1px solid #4d90fe;outline:rgba(0,0,0,0) 0}.ndfHFb-c4YZDc-Sx9Kwc-c6xFrd .ndfHFb-c4YZDc-ldDVFe-JIbuQc[disabled]{-moz-box-shadow:none;box-shadow:none;background:#4d90fe;color:#fff;filter:alpha(opacity=50);opacity:.5}.ndfHFb-c4YZDc-Sx9Kwc-TD02Lb{position:absolute;visibility:hidden}.VIpgJd-TUo6Hb,.XKSfm-Sx9Kwc{-moz-box-shadow:0 4px 16px rgba(0,0,0,.2);box-shadow:0 4px 16px rgba(0,0,0,.2);background:#fff;background-clip:padding-box;border:1px solid #acacac;border:1px solid rgba(0,0,0,.333);outline:0;position:absolute}.VIpgJd-TUo6Hb-xJ5Hnf,.XKSfm-Sx9Kwc-xJ5Hnf{background:#fff;left:0;position:absolute;top:0}div.VIpgJd-TUo6Hb-xJ5Hnf,div.XKSfm-Sx9Kwc-xJ5Hnf{filter:alpha(opacity=75);opacity:.75}.XKSfm-Sx9Kwc{color:#000;padding:30px 42px}.XKSfm-Sx9Kwc-r4nke{background-color:#fff;color:#000;cursor:default;font-size:16px;font-weight:normal;line-height:24px;margin:0 0 16px}.XKSfm-Sx9Kwc-r4nke-TvD9Pc{height:11px;opacity:.7;padding:17px;position:absolute;right:0;top:0;width:11px}.XKSfm-Sx9Kwc-r4nke-TvD9Pc:after{content:"";background:url(//ssl.gstatic.com/ui/v1/dialog/close-x.png);position:absolute;height:11px;width:11px;right:17px}.XKSfm-Sx9Kwc-r4nke-TvD9Pc:hover{opacity:1}.XKSfm-Sx9Kwc-bN97Pc{background-color:#fff;line-height:1.4em;word-wrap:break-word}.XKSfm-Sx9Kwc-c6xFrd{margin-top:16px}.XKSfm-Sx9Kwc-c6xFrd button{-moz-border-radius:2px;border-radius:2px;background-color:#f5f5f5;background-image:-moz-linear-gradient(top,#f5f5f5,#f1f1f1);background-image:linear-gradient(top,#f5f5f5,#f1f1f1);border:1px solid #dcdcdc;border:1px solid rgba(0,0,0,.1);color:#444;cursor:default;font-family:inherit;font-size:11px;font-weight:bold;height:29px;line-height:27px;margin:0 16px 0 0;min-width:72px;outline:0;padding:0 8px}.XKSfm-Sx9Kwc-c6xFrd button:hover{-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1);background-color:#f8f8f8;background-image:-moz-linear-gradient(top,#f8f8f8,#f1f1f1);background-image:linear-gradient(top,#f8f8f8,#f1f1f1);border:1px solid #c6c6c6;color:#333}.XKSfm-Sx9Kwc-c6xFrd button:active{-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1);background-color:#f8f8f8;background-image:-moz-linear-gradient(top,#f8f8f8,#f1f1f1);background-image:linear-gradient(top,#f8f8f8,#f1f1f1);border:1px solid #c6c6c6;color:#333;-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.1);box-shadow:inset 0 1px 2px rgba(0,0,0,.1)}.XKSfm-Sx9Kwc-c6xFrd button:focus{border:1px solid #4d90fe}.XKSfm-Sx9Kwc-c6xFrd button[disabled]{-moz-box-shadow:none;box-shadow:none;background:#fff;background-image:none;border:1px solid #f3f3f3;border:1px solid rgba(0,0,0,.05);color:#b8b8b8}.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc{background-color:#4d90fe;background-image:-moz-linear-gradient(top,#4d90fe,#4787ed);background-image:linear-gradient(top,#4d90fe,#4787ed);border:1px solid #3079ed;color:#fff}.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:hover{background-color:#357ae8;background-image:-moz-linear-gradient(top,#4d90fe,#357ae8);background-image:linear-gradient(top,#4d90fe,#357ae8);border:1px solid #2f5bb7;color:#fff}.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:active{background-color:#357ae8;background-image:-moz-linear-gradient(top,#4d90fe,#357ae8);background-image:linear-gradient(top,#4d90fe,#357ae8);border:1px solid #2f5bb7;color:#fff;-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.3);box-shadow:inset 0 1px 2px rgba(0,0,0,.3)}.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:focus{-moz-box-shadow:inset 0 0 0 1px #fff;box-shadow:inset 0 0 0 1px #fff;border:1px solid #fff;border:rgba(0,0,0,0) solid 1px;outline:1px solid #4d90fe;outline:rgba(0,0,0,0) 0}.XKSfm-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc[disabled]{-moz-box-shadow:none;box-shadow:none;background:#4d90fe;color:#fff;filter:alpha(opacity=50);opacity:.5}.tk3N6e-O0r3Gd,.tk3N6e-McfNlf,.tk3N6e-ostUZ{width:512px}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;align-items:flex-start;padding-bottom:16px;outline:none;position:absolute;width:384px;height:auto;background:#fff;-moz-box-shadow:0 1px 2px rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);box-shadow:0 1px 2px rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);-moz-border-radius:8px;border-radius:8px;z-index:1195}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-bN97Pc{max-width:100%}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-xJ5Hnf{background-color:#000;height:100%;left:0;position:fixed;top:0;width:100%;z-index:1194}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-r4nke{margin:0 auto}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -64px;width:24px;height:24px;margin:18px auto 10px;transform:scale(1.3)}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-r4nke-fmcmS{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;letter-spacing:0;line-height:1.75rem;color:#202124}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-C7uZwb-bN97Pc{letter-spacing:.01428571em;font-family:Roboto,Arial,sans-serif;font-size:.875rem;font-weight:400;line-height:1.25rem;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;height:100px;flex-direction:column;margin:16px 24px 20px;justify-content:space-around}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-hSRGPd{color:#5f6368;overflow:hidden;text-overflow:ellipsis}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-Ne3sFf{color:#202124}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-KY1xSc-z5C9Gb{font-weight:100;margin:0 5px;position:relative;top:-2px}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-c6xFrd{margin-left:auto;margin-right:24px}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-ssJRIf-LgbsSe:hover,.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-K4efff-LgbsSe:hover{cursor:pointer}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-ssJRIf-LgbsSe{font-family:"Google Sans",Roboto,arial,sans-serif;text-align:center;min-width:70px;background:#f9ab00;-moz-border-radius:5px;border-radius:5px;font-size:14px;padding:8px 24px;border-style:none;outline:none}.ndfHFb-c4YZDc-uWtm3-GMvhG-Sx9Kwc-K4efff-LgbsSe{font-family:"Google Sans",Roboto,arial,sans-serif;margin:0 16px;text-align:center;min-width:70px;font-size:14px;padding:7px 0;border-style:none;background:#fff;outline:none}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{color:rgba(255,255,255,0.87);font-size:11px;font-weight:bold;text-align:center;text-shadow:0 1px 0 rgba(0,0,0,.8);vertical-align:middle;height:27px;line-height:27px;margin-right:2px;min-width:50px;padding:10px 0}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{text-shadow:none}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{-moz-border-radius:2px;border-radius:2px;height:24px;line-height:24px;margin:0;padding:8px;min-width:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{-moz-border-radius:100px;border-radius:100px}.ndfHFb-c4YZDc-AHmuwe-Hr88gd-qnnXGd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe{border-color:#575757}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-AHmuwe-Hr88gd-qnnXGd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe{background-color:rgba(196,199,197,.12)}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me{color:rgba(255,255,255,0.47);text-shadow:none}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{color:rgba(255,255,255,1);background-color:#232323;background-image:-moz-linear-gradient(top,#333,#222);background-image:linear-gradient(top,#333,#222)}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:#838383;background-image:none}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd{-moz-box-shadow:inset 0 1px 6px rgba(0,0,0,.8);box-shadow:inset 0 1px 6px rgba(0,0,0,.8)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-LgbsSe-auswjd{-moz-box-shadow:none;box-shadow:none;background-color:rgba(255,255,255,.35)}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-LgbsSe-auswjd{background-color:rgba(196,199,197,.12)}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe{background-color:rgba(35,35,35,.6);border-bottom:3px solid #4d90fe;padding-bottom:7px}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe{background-color:#6d6e71;border-bottom-color:#58595b}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:#838383}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{-moz-transition:background-color 0.1s,opacity 0.1s;transition:background-color 0.1s,opacity 0.1s}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:rgba(255,255,255,.25);background-image:none}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:rgba(196,199,197,.08)}.ndfHFb-c4YZDc-LgbsSe-IwzHHe .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe,.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe{background-color:rgba(255,255,255,.1);border-bottom-color:#c1d9ff}.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd,.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-auswjd{-moz-box-shadow:inset 0 1px 6px rgba(0,0,0,.4);box-shadow:inset 0 1px 6px rgba(0,0,0,.4)}.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE,.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE,.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe,.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe{background:#609cfd;outline:0}.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd .ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe{background:#1f59c0}.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd{display:inline-block;margin:6px 0}.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-to915-LgbsSe{background-color:#3f76d9}.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background:#407ff1}.ndfHFb-c4YZDc-Wrql6b-gvZm2b-c6xFrd .ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-JbbQac.ndfHFb-c4YZDc-to915-LgbsSe{margin-right:1px;min-width:35px;width:35px;padding:4px 0;margin-left:5px}.ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-JbbQac .ndfHFb-c4YZDc-Bz112c{background-position:0 0;width:25px;height:25px;padding:3px 10px;margin-left:4px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-JbbQac .ndfHFb-c4YZDc-Bz112c{background-position:0 -1528px}.ndfHFb-c4YZDc-Wrql6b-gvZm2b-LgbsSe-V67aGc{font-size:13px;text-transform:uppercase;text-shadow:none;color:white;display:inline-block;padding-left:3px}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-Wrql6b-gvZm2b-xl07Ob-LgbsSe{padding:4px 10px;margin-right:5px}.ndfHFb-c4YZDc-Wrql6b-gvZm2b-xl07Ob-LgbsSe .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo{margin-left:5px}.ndfHFb-c4YZDc .ndfHFb-aZ2wEe{display:none;height:100%;width:100%}.ndfHFb-c4YZDc .ndfHFb-vyDMJf-aZ2wEe{height:21px;margin-left:-10.5px;top:0;width:21px}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-vyDMJf-aZ2wEe{height:24px;margin-left:-12px;width:24px}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb{display:inline-block}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb{z-index:1;display:none}.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c{background-repeat:no-repeat;filter:alpha(opacity=87);opacity:0.87;margin-left:auto;margin-right:auto;margin-top:3px;height:21px;width:21px}.ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c{background-repeat:no-repeat;filter:alpha(opacity=87);opacity:0.87;margin-left:auto;margin-right:auto;height:21px}.ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c{background-repeat:no-repeat;filter:alpha(opacity=87);opacity:0.87;margin-left:auto;margin-right:auto;margin-top:3px;height:21px;width:21px}.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c,.ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c,.ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c{background-repeat:no-repeat;filter:alpha(opacity=87);opacity:0.87;margin-left:auto;margin-right:auto;margin-top:2px;height:24px;width:24px}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg')!important}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/v-spinner_dark.gif')!important}.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c{background-position:0 -240px}.ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c{background-position:0 -600px}.ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c{background-position:0 -400px}.ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c{background-position:0 -1920px}.ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c{margin-top:4px;width:19px}.ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c{background-position:0 -2360px}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited){margin-top:2px;height:24px;width:24px;background-image:none!important;filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c .ndfHFb-aZ2wEe{display:block}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-mJSDk-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-w37qKe-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg')!important}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-mJSDk-wcotoc-ndfHFb-Bz112c{background-position:0 -1816px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c{background-position:0 -1448px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c{background-position:0 -896px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c{background-position:0 -1568px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-w37qKe-Bz112c{background-position:0 -448px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c{background-position:0 -328px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c{background-position:0 -2464px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-mJSDk-wcotoc-ndfHFb-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-mvmHBc-wcotoc-ndfHFb-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-x5cW0b-wcotoc-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-w37qKe-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-ndfHFb-w37qKe-Bz112c{filter:alpha(opacity=100);opacity:1;margin-top:0;height:24px;width:24px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c{filter:alpha(opacity=100);opacity:1;margin:2.5px;width:19px;height:19px}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-KJlZme-wcotoc-ndfHFb-Bz112c:not([onclick]):not(:link):not(:visited){margin:0;height:24px;width:24px}.ndfHFb-c4YZDc-Sx9Kwc.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc{padding:0}.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-r4nke{border-bottom:1px solid #acacac;font-family:arial,sans-serif;padding:15px 12px}.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde{background-color:#f3f3f3;height:100%;position:relative;width:100%}.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde .ndfHFb-c4YZDc-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde-k4Qmrd{text-align:center;width:100%;position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-DWWcKd-ZpdDCc-ge6pde-RJLb9c{background-image:url('//ssl.gstatic.com/ui/v1/activityindicator/loading_bg_f5.gif');background-repeat:no-repeat;display:inline-block;height:19px;position:relative;top:3px;width:19px}.ndfHFb-c4YZDc-y0R6E-DWWcKd-b3rLgd{display:inline-block;vertical-align:middle}.ndfHFb-c4YZDc-y0R6E-DWWcKd-Bz112c{display:inline-block;height:12px;width:12px}.ndfHFb-c4YZDc-y0R6E-DWWcKd-Ne3sFf{display:inline-block;padding-left:16px;vertical-align:top}.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-xJ5Hnf{background-color:#202124;left:0;position:absolute;top:0;z-index:1194}.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc{background-color:#fff;-moz-border-radius:8px;border-radius:8px;font-family:"Google Sans",Roboto,arial,sans-serif;padding:20px;position:absolute;width:450px;z-index:1195}.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-c6xFrd{float:right;margin-top:20px}.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-LgbsSe{background:#fff;border-color:#bdc1c6;-moz-border-radius:4px;border-radius:4px;border-style:solid;border-width:1px;color:#1a73e8;cursor:pointer;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;line-height:2;margin-left:5px;padding:0 20px}.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-zTETae{background:#1a73e8;color:#fff}.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-r4nke-fmcmS{font-size:22px}.ndfHFb-c4YZDc-RvPyde-S9gUrf-Sx9Kwc-bN97Pc{color:#5f6368;font-size:14px;margin:10px 0}.ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf{align-items:center;background:#e8f0fe;color:#202124;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;font-family:"Google Sans",Roboto,arial,sans-serif;height:48px;width:100%}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf{background:#7cacf8}.ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf.ndfHFb-c4YZDc-MqcBrc-ORHb-L6cTce,.ndfHFb-c4YZDc-MqcBrc-ORHb-c6xFrd.ndfHFb-c4YZDc-MqcBrc-ORHb-L6cTce,.ndfHFb-c4YZDc-MqcBrc-ORHb-L6cTce{display:none}.ndfHFb-c4YZDc-MqcBrc-ORHb-c6xFrd{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:1;flex-grow:1;float:right;justify-content:flex-end}.ndfHFb-c4YZDc-MqcBrc-ORHb-Bz112c{background-position:0 -2544px;height:24px;margin:0 16px;width:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-Bz112c{background-position:0 -3634px}.ndfHFb-c4YZDc-MqcBrc-ORHb-Vkfede-Ne3sFf{margin-left:16px;font-size:14px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-Vkfede-Ne3sFf{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-MqcBrc-ORHb-jOfkMb{font-size:16px;font-weight:500}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-jOfkMb{font:var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-title-medium-spacing,0.00625em)}.ndfHFb-c4YZDc-MqcBrc-ORHb-IYtByb-LgbsSe-Bz112c{background-position:0 -1160px;height:24px;width:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-IYtByb-LgbsSe-Bz112c{background-position:0 -3570px;height:20px;width:24px}.ndfHFb-c4YZDc-MqcBrc-ORHb-IYtByb-LgbsSe-sM5MNb{margin:0 16px}.ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe:hover,.ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe:hover{cursor:pointer}.ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe{margin:0 12px;text-align:center;min-width:70px;background:#1a73e8;-moz-border-radius:5px;border-radius:5px;font-size:14px;font-weight:500;padding:7px 0;color:#fff}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe{margin:0 12px;color:#202124;background:none;font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em)}.ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe:hover{background:#2b7de9}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-ssJRIf-LgbsSe:hover{background:none}.ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe{margin:0 5px;text-align:center;min-width:70px;color:#1a73e8;font-size:14px;font-weight:500;padding:7px 0}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe{margin:0 12px;color:#202124;background:none;font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em)}.ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe:hover{background:#f8fbff}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MqcBrc-ORHb-K4efff-LgbsSe:hover{background:none}.ndfHFb-c4YZDc-rovI0b{color:#fff;font-size:13px;font-weight:normal;text-align:left;text-shadow:0px 2px 1px rgba(0,0,0,.1);white-space:nowrap}.ndfHFb-c4YZDc-rovI0b-r4nke{line-height:30px;margin-bottom:10px;text-align:center}.ndfHFb-c4YZDc-rovI0b-bN97Pc{overflow-x:hidden;overflow-y:auto;border-top:1px solid #696868;border-bottom:1px solid #696868;min-height:55px}.ndfHFb-c4YZDc-rovI0b-bN97Pc.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb{min-height:0!important}.ndfHFb-c4YZDc-rovI0b-LS81yb{padding-bottom:10px}.ndfHFb-c4YZDc-rovI0b-LS81yb-Ud7fr{border-bottom:none;color:#cdcdcd;font-size:13px;font-weight:normal;line-height:25px;padding:0}.ndfHFb-c4YZDc-rovI0b-IyROMc-rymPhb{margin-left:100px}.ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b{cursor:pointer;display:block;padding:6px 15px 6px 0;border:none}.ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b.ndfHFb-c4YZDc-w5vlXd{border:none}.ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b:hover{background-color:#444;border-color:#444;border-style:dotted;border-width:1px 0;padding:5px 15px 5px 0}.ndfHFb-c4YZDc-rovI0b-ljLd3-IyROMc .ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b{font-weight:bold}.ndfHFb-c4YZDc-rovI0b-UEIKff-IyROMc .ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b,.ndfHFb-c4YZDc-rovI0b-MVH0Ye-IyROMc .ndfHFb-c4YZDc-rovI0b-DWWcKd-ibnC6b{font-weight:normal}.ndfHFb-c4YZDc-rovI0b-DWWcKd-Bz112c{display:inline-block;height:16px;margin-left:5px;vertical-align:middle;width:16px}.ndfHFb-c4YZDc-rovI0b-DWWcKd-V1ur5d{display:inline-block;line-height:16px;margin-left:20px}.ndfHFb-c4YZDc-JqEhuc-s2gQvd{bottom:0;overflow:auto;position:absolute}.ndfHFb-c4YZDc-JqEhuc{background-color:#fff;border:20px solid transparent;-moz-border-radius:20px;border-radius:20px;color:#000;font-size:14px;position:absolute;word-wrap:break-word;-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35)}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-JqEhuc{border:none;-moz-border-radius:0;border-radius:0;border-top:10px solid transparent;-moz-box-shadow:none;box-shadow:none}.ndfHFb-c4YZDc-JqEhuc-bN97Pc,.ndfHFb-c4YZDc-JqEhuc-tJHJj{margin-left:20px;margin-right:20px;right:0;left:0}.ndfHFb-c4YZDc-JqEhuc-n5VRYe{background-color:none;background-image:-moz-linear-gradient(rgba(0,0,0,.2),transparent);background-image:linear-gradient(rgba(0,0,0,.2),transparent);height:8px;left:20px;position:absolute;right:20px;z-index:1}.ndfHFb-c4YZDc-JqEhuc-r4nke{display:inline-block;font-size:30px;margin-right:10px;margin-left:10px;max-width:85%;filter:alpha(opacity=60);opacity:.6;overflow:hidden;padding-bottom:10px;text-overflow:ellipsis;vertical-align:middle}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-r4nke{line-height:50px;padding-bottom:0}.ndfHFb-c4YZDc-JqEhuc-r4nke-tJHJj{border-bottom:1px solid #cececf}.ndfHFb-c4YZDc-JqEhuc-r4nke-oKdM2c{filter:alpha(opacity=60);opacity:.6;font-size:10px;display:block;overflow:hidden;white-space:nowrap}.ndfHFb-c4YZDc-JqEhuc-NnAfwf{display:inline-block;font-size:16px;filter:alpha(opacity=60);opacity:.6;vertical-align:middle}.ndfHFb-c4YZDc-JqEhuc-oKdM2c,.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c{border-bottom:1px solid #cececf;display:block;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c.ndfHFb-c4YZDc-LgbsSe{display:block}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-tJHJj .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c{height:50px}.ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe,.ndfHFb-c4YZDc-JqEhuc-PlOyMe-Bz112c.ndfHFb-c4YZDc-LgbsSe,.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-JqEhuc-oKdM2c,.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c{cursor:pointer}.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-JqEhuc-oKdM2c,.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c,.ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe:hover,.ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe:active,.ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe{background-color:#ddd}.ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-oKdM2c,.ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-bMcfAe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-oKdM2c,.ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c,.ndfHFb-c4YZDc-JqEhuc-bN97Pc .ndfHFb-c4YZDc-bMcfAe-ZmdkE.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c{background-color:#e8f0fe;color:#185abc}.ndfHFb-c4YZDc-JqEhuc-oKdM2c-Bz112c{background-size:contain;display:inline-block;height:16px;width:16px;margin-left:10px;margin-right:10px;position:relative;top:3px}.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-Bz112c{background-size:contain;display:inline-block;height:16px;width:16px;margin-left:3%;margin-right:3%;position:relative;top:10px}.ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c{background-position:0 -1840px;height:21px;width:21px;left:-5px;top:8px;position:absolute}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c{background-position:0 -1080px}.ndfHFb-c4YZDc-JqEhuc-oKdM2c-V1ur5d{display:inline;line-height:38px}.ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb{float:left}.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d,.ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd,.ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe{display:inline-block;line-height:38px;overflow:hidden;text-overflow:ellipsis}.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d{width:50%}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d{font-size:12px}.ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd{width:22%;filter:alpha(opacity=60);opacity:.6}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd{font-size:12px;opacity:1}.ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe{width:13%;filter:alpha(opacity=60);opacity:.6}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe{font-size:12px;opacity:1}.ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c:after{content:"";display:table;clear:both}.ndfHFb-c4YZDc-kODWGd{position:absolute}.ndfHFb-c4YZDc-kODWGd-nK2kYb{-moz-user-select:none;-moz-border-radius:5px;border-radius:5px;background-color:rgba(20,20,20,.8);position:absolute;height:100%;width:100%;-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35)}.ndfHFb-c4YZDc-kODWGd-NziyQe-LgbsSe{position:absolute;top:2px;left:10px;right:auto}.ndfHFb-c4YZDc-kODWGd-HvfI2b-Bz112c{height:28px;width:26px}.ndfHFb-c4YZDc-kODWGd-NziyQe-Bz112c{height:28px;width:26px;background-position:0 -1120px}.ndfHFb-c4YZDc-kODWGd-HvfI2b-Bz112c{background-position:0 -120px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-NziyQe-Bz112c{background-position:0 -3386px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-HvfI2b-Bz112c{background-position:0 -2344px}.ndfHFb-c4YZDc-kODWGd-bVEB4e{border:1px solid #b3b3b3;background-color:#0a0a0a;display:table-cell;pointer-events:auto;text-align:center;vertical-align:middle}.ndfHFb-c4YZDc-kODWGd-LgbsSe{-moz-border-radius:0;border-radius:0;-moz-transition:all .218s;transition:all .218s;background-color:#f3f3f3;border:1px solid rgba(0,0,0,.1);color:#444;font-weight:bold;font-size:11px;height:27px;line-height:27px;margin:6px;min-width:54px;padding:0 8px;text-align:center}.ndfHFb-c4YZDc-kODWGd-LgbsSe:hover{background-color:#d8d8d8;border:1px solid #c6c6c6;color:#222;-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1)}.ndfHFb-c4YZDc-kODWGd-nK2kYb .ndfHFb-c4YZDc-SxecR{padding-left:0px!important;padding-right:2px!important}.ndfHFb-c4YZDc-kODWGd-nK2kYb .ndfHFb-c4YZDc-SxecR-skjTt-MFS4be{border-bottom-left-radius:8px!important;border-top-left-radius:8px!important;border-bottom-right-radius:0px!important;border-top-right-radius:0px!important;padding-left:0px!important;padding-right:3px!important}.ndfHFb-c4YZDc-TL3Ynd-V67aGc-haAclf{display:inline-block}.ndfHFb-c4YZDc-TL3Ynd-V67aGc{cursor:pointer;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;margin-left:16px}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-haAclf{display:block;position:absolute;white-space:normal}.ndfHFb-c4YZDc-Btuy5e-Rgw69b{margin-left:16px;top:11px}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-L6cTce{visibility:hidden}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-TvD9Pc-LgbsSe{-moz-border-radius:24px;border-radius:24px;height:24px;padding:12px;width:24px;z-index:1194}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-TvD9Pc-LgbsSe:hover{background:#f1f3f4}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-TvD9Pc-LgbsSe:active{background:#dadce0}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-fmcmS-LgbsSe{align-items:center;-moz-border-radius:2px;border-radius:2px;color:#1a73e8;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;font-size:14px;height:36px;letter-spacing:.15px;margin:6px 0;min-width:60px;outline:1px solid transparent;padding:0 15px;z-index:1194}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-fmcmS-LgbsSe:hover{background:#e8f0fe}.ndfHFb-c4YZDc-Btuy5e-Rgw69b-fmcmS-LgbsSe:active{background:#d2e3fc}.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar{height:12px;overflow:visible;width:12px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar{width:16px}.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-button{height:0;width:0}.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-corner{background:transparent}.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-track{background-color:transparent;-moz-box-shadow:none!important;box-shadow:none!important;border:none}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-track{background-color:rgba(255,255,255,.1)}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-track{background:transparent}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-thumb{background-color:rgba(255,255,255,.9)}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-track{background-color:rgba(0,0,0,.1)}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-sn54Q::-webkit-scrollbar-thumb{background-color:rgba(0,0,0,.6)}.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb{background-color:#4c4c4c;background-clip:padding-box;border-style:solid;border-color:transparent;border-width:0 1px 0 0;-moz-box-shadow:inset 1px 1px 0 #676767,inset 0 -1px 0 #676767;box-shadow:inset 1px 1px 0 #676767,inset 0 -1px 0 #676767;min-height:75px;padding:100px 0 0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb{background-color:rgba(255,255,255,.75);-moz-border-radius:1px;border-radius:1px;border-width:0;-moz-box-shadow:none;box-shadow:none;min-height:56px;padding:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb{background-color:var(--dt-outline-variant,#dadce0);-moz-border-radius:100px;border-radius:100px;border:solid 4px transparent;background-clip:padding-box}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb{background-color:rgba(0,0,0,.5)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-to915::-webkit-scrollbar-thumb{background-color:#4c4c4c}.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb:hover{background-color:#9f9f9f;-moz-box-shadow:inset 1px 1px 0 #ccc;box-shadow:inset 1px 1px 0 #ccc}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb:hover{background-color:rgba(255,255,255,.9);-moz-box-shadow:none;box-shadow:none}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-thumb:hover{background-color:var(--dt-outline-variant,#dadce0)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-s2gQvd.ndfHFb-c4YZDc-s2gQvd-to915::-webkit-scrollbar-thumb:hover{background-color:#9f9f9f}.ndfHFb-c4YZDc-s2gQvd{scrollbar-face-color:#666;scrollbar-track-color:#2e2e2e;scrollbar-arrow-color:#666;scrollbar-shadow-color:#717171}.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar{display:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-cYSp0e-s2gQvd.ndfHFb-c4YZDc-s2gQvd::-webkit-scrollbar-track-piece:start{margin-top:64px}.ndfHFb-c4YZDc-MqcBrc-ORHb-haAclf.ndfHFb-c4YZDc-ORHb-L6cTce,.ndfHFb-c4YZDc-uWtm3-ORHb.ndfHFb-c4YZDc-ORHb-L6cTce,.ndfHFb-c4YZDc-ORHb-L6cTce{display:none}.ndfHFb-c4YZDc-uWtm3-ORHb{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;background-color:#f9ab00;-moz-border-radius:0;border-radius:0;color:#202124;height:3rem;position:relative;top:0;width:100%;z-index:3}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb{background:#ffdf99}.ndfHFb-c4YZDc-uWtm3-ORHb-bN97Pc{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;justify-content:space-between;width:100%}.ndfHFb-c4YZDc-uWtm3-ORHb-Ne3sFf{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-Ne3sFf{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-uWtm3-ORHb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -1240px;height:24px;margin:0 25px;width:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-Bz112c{margin:0 16px}.ndfHFb-c4YZDc-uWtm3-ORHb-LQLjdd{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;align-items:center;margin:8px 0;-moz-box-ordinal-group:0;order:0}.ndfHFb-c4YZDc-uWtm3-ORHb-IYtByb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3570px;height:20px;margin:0 25px;width:20px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-IYtByb-Bz112c{margin:0 16px;height:20px;width:24px}.ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe,.ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe{align-self:center;color:#202124;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px;padding:0 8px;text-align:center;text-decoration:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe{font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em);padding:0 12px}.ndfHFb-c4YZDc-uWtm3-ORHb-GrFcDd-ShBeI-LgbsSe:hover,.ndfHFb-c4YZDc-uWtm3-ORHb-KY1xSc-z5C9Gb-LgbsSe:hover{cursor:pointer}.ndfHFb-c4YZDc-wvGCSb-gkA7Yd{right:-50px;position:absolute;width:49px;top:0;z-index:3}.ndfHFb-c4YZDc-RDNXzf-L6cTce .ndfHFb-c4YZDc-wvGCSb-gkA7Yd{display:none}.ndfHFb-c4YZDc-VCkuzd{min-height:190px;width:500px;bottom:10px;position:absolute;right:10px;z-index:10;-moz-box-shadow:0 0 20px rgba(0,0,0,.8);box-shadow:0 0 20px rgba(0,0,0,.8);background-color:#fff;padding:10px}.ndfHFb-c4YZDc-VCkuzd::after{content:"";height:0;width:0;bottom:-18px;right:5%;position:absolute;border-top:18px solid #fff;border-left:15px solid transparent;border-right:15px solid transparent}.ndfHFb-c4YZDc-eLiUMc-Tswv1b-haAclf{margin-bottom:6px;margin-right:6px;vertical-align:top}.ndfHFb-c4YZDc-eLiUMc-Tswv1b{color:#777;font-size:8px}.ndfHFb-c4YZDc-eLiUMc-Tswv1b-haAclf.ndfHFb-c4YZDc-eLiUMc-Tswv1b{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;position:absolute;right:0;bottom:0;z-index:1293}.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd{-moz-border-radius:2px;border-radius:2px;border:0 solid;-moz-box-shadow:0px 2px 4px rgba(0,0,0,.2);box-shadow:0px 2px 4px rgba(0,0,0,.2);display:none;height:0;visibility:hidden;font-size:11px;overflow:hidden;padding:0;text-align:center;-moz-transition:all 0 linear 1s,opacity 1s;transition:all 0 linear 1s,opacity 1s;background-color:#f9edbe;border-color:#f0c36d;color:#333}.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-TSZdd{-moz-transition:opacity 0.218s;transition:opacity 0.218s;border-width:1px;display:inline-block;height:auto;max-width:90%;padding:6px 16px;text-overflow:ellipsis;visibility:visible}.ndfHFb-c4YZDc-X3SwIb.ndfHFb-c4YZDc-b3rLgd-haAclf{height:0;position:absolute;text-align:center;top:50px;width:100%;z-index:4}.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd{padding-left:6px}.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd,.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-hSRGPd,.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited,.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-hSRGPd:visited{color:#00f;cursor:pointer;text-decoration:none}.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover,.ndfHFb-c4YZDc-X3SwIb .ndfHFb-c4YZDc-b3rLgd-hSRGPd:hover{text-decoration:underline}.ndfHFb-c4YZDc-LgbsSe{cursor:default}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe{cursor:pointer;display:inline-block}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-OWB6Me{cursor:default}.ndfHFb-c4YZDc-jNm5if-Hn6s1b{background:rgba(66,133,244,.9);border-color:transparent;-moz-border-radius:50%;border-radius:50%;border-style:solid;border-width:30px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;height:320px;justify-content:center;position:absolute;right:-25px;top:-72px;white-space:normal;width:320px;z-index:10}.ndfHFb-c4YZDc-jNm5if-Hn6s1b-bBybbf{height:100%;width:100%;position:relative;z-index:10}.ndfHFb-c4YZDc-jNm5if-Hn6s1b .ndfHFb-c4YZDc-jNm5if-Hn6s1b-tJHJj{font-size:20px;font-weight:normal;line-height:24px}.ndfHFb-c4YZDc-jNm5if-Hn6s1b .ndfHFb-c4YZDc-jNm5if-Hn6s1b-Ne3sFf{font-size:14px;line-height:24px}.ndfHFb-c4YZDc-jNm5if-Hn6s1b-LgbsSe{position:absolute}.ndfHFb-c4YZDc-jNm5if-Hn6s1b-LgbsSe-Bz112c{background-position:0 -1632px;height:24px;left:32px;opacity:.6;position:relative;top:34px;width:24px}.ndfHFb-c4YZDc-jNm5if-Hn6s1b-LgbsSe-LkdAo{background:white;-moz-border-radius:50%;border-radius:50%;height:88px;left:-32px;position:absolute;top:-34px;width:88px}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b{animation:expandCallout .6s;-moz-border-radius:50%;border-radius:50%;color:white;justify-content:center;line-height:24px;position:absolute;transition:all ease-out;white-space:normal}@keyframes expandCallout{0%{transform:scale(0,0)}to{transform:scale(1,1)}}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b-bBybbf{height:100%;position:relative;width:100%;z-index:2}.UMrnmb-v3pZbf .ndfHFb-c4YZDc-FNFY6c-Hn6s1b{-moz-box-shadow:0 100px 0 250px rgba(17,109,231,.96);box-shadow:0 100px 0 250px rgba(17,109,231,.96)}.UMrnmb-nllRtd .ndfHFb-c4YZDc-FNFY6c-Hn6s1b{-moz-box-shadow:0 100px 0 250px rgba(21,138,54,.96);box-shadow:0 100px 0 250px rgba(21,138,54,.96)}.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-FNFY6c-Hn6s1b{-moz-box-shadow:0 100px 0 250px rgba(249,168,0,.96);box-shadow:0 100px 0 250px rgba(249,168,0,.96);color:black}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-bN97Pc{background-color:rgba(0,0,0,.005);border:1px solid transparent;padding:0 30px 30px 30px;width:400px}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-tJHJj{font-size:20px;font-weight:normal;margin-bottom:10px}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-Ne3sFf{font-size:14px}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-KY1xSc-z5C9Gb{color:white;display:inline-block;font-size:14px;font-weight:bold;margin-left:10px;text-decoration:none}.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-KY1xSc-z5C9Gb{color:black}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-c6xFrd{font-size:14px;font-weight:bold}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-iDjqhe-Hnhb3b-WtFGnf{border:1px solid transparent;display:inline-block}.ndfHFb-c4YZDc-FNFY6c-Hn6s1b .ndfHFb-c4YZDc-FNFY6c-Hn6s1b-F2rEXb{border:1px solid transparent;display:inline-block;margin-left:40px;opacity:.75}.UMrnmb-v3pZbf .ndfHFb-c4YZDc-G0brRe-Hn6s1b{background-color:rgba(17,109,231,.96)}.UMrnmb-nllRtd .ndfHFb-c4YZDc-G0brRe-Hn6s1b{background-color:rgba(21,138,54,.96)}.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-G0brRe-Hn6s1b{background-color:rgba(249,168,0,.96);color:black}.ndfHFb-c4YZDc-G0brRe-Hn6s1b{-moz-border-radius:4px 0 0 4px;border-radius:4px 0 0 4px;height:40px;margin:0 auto;position:absolute;right:0;top:56px}.ndfHFb-c4YZDc-G0brRe-Hn6s1b-Ne3sFf{float:left;font-size:14px;line-height:40px;margin-bottom:0;margin-top:0;padding:0 32px 0 24px}.ndfHFb-c4YZDc-G0brRe-Hn6s1b-scrj1b-G0brRe{color:white;font-size:14px;font-weight:bold;line-height:40px;margin-bottom:0;margin-top:0}.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-G0brRe-Hn6s1b-scrj1b-G0brRe{color:black}.UMrnmb-gS7Ybc .ndfHFb-c4YZDc-G0brRe-Hn6s1b-TvD9Pc{background-position:0 -1120px}.ndfHFb-c4YZDc-G0brRe-Hn6s1b-TvD9Pc{background-position:0 -3178px;float:right;height:20px;margin-left:32px;margin-right:24px;margin-top:8px;opacity:.5;width:20px}.ndfHFb-c4YZDc-K9a4Re-nKQ6qf{position:absolute;top:0;bottom:0;width:100%;-moz-user-select:none}.ndfHFb-c4YZDc-K9a4Re-ge6pde-Ne3sFf{position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-oKVyEf{-moz-user-select:text}.ndfHFb-c4YZDc-MZArnb-b0t70b{-moz-box-sizing:border-box;box-sizing:border-box;-moz-box-shadow:inset 0 0 10px #000;box-shadow:inset 0 0 10px #000;background-color:#242223;bottom:0;position:fixed;right:0;top:47px;width:400px;z-index:1}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b{-moz-box-shadow:none;box-shadow:none;background-color:#323232;width:344px;top:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b{background:none;padding:0 16px 16px 0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b-haAclf{background:var(--dt-surface,#fff);-moz-border-radius:24px;border-radius:24px;height:100%;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-MZArnb-b0t70b{z-index:4}.ndfHFb-c4YZDc-MZArnb-b0t70b-L6cTce{display:none}.ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c{display:block;margin-left:auto;margin-right:auto}.ndfHFb-c4YZDc-MZArnb-tJHJj{-moz-box-sizing:border-box;box-sizing:border-box;font-family:Roboto,arial,sans-serif;font-size:14px;text-transform:uppercase}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-tJHJj{-moz-box-shadow:0 2px 2px rgba(0,0,0,.3);box-shadow:0 2px 2px rgba(0,0,0,.3);font-family:"Google Sans",Roboto,arial,sans-serif;font-size:16px;text-transform:none}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-tJHJj{-moz-box-shadow:none;box-shadow:none;border-bottom:solid 2px var(--dt-outline-variant,#dadce0)}.ndfHFb-c4YZDc-MZArnb-bN97Pc{bottom:0;left:0;margin:5px 0;overflow-y:auto;position:absolute;right:0;top:50px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-MZArnb-bN97Pc{position:static;top:0;margin:5px 0 15px 0}.ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e{-moz-box-sizing:border-box;box-sizing:border-box;color:#c0bebe;cursor:pointer;display:inline-block;height:50px;line-height:50px;margin:0 16px 0;padding:4px 2px 0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e{height:56px;line-height:56px}.ndfHFb-c4YZDc-MZArnb-cXCLoc{border-bottom:1px solid #ccc;margin:0 15px 0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-cXCLoc{border-bottom:none;display:inline-block;margin:0}.ndfHFb-c4YZDc-MZArnb-AznF2e-gk6SMd.ndfHFb-c4YZDc-MZArnb-AznF2e-uDEFge{border-bottom:3px solid #4d90fe}.ndfHFb-c4YZDc-MZArnb-AznF2e:hover.ndfHFb-c4YZDc-MZArnb-AznF2e-uDEFge{border-bottom:3px solid #646464}.ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e:hover{margin:0 18px 0;padding:4px 0 0}.ndfHFb-c4YZDc-MZArnb-tJHJj .ndfHFb-c4YZDc-MZArnb-AznF2e.ndfHFb-c4YZDc-MZArnb-AznF2e-gk6SMd{color:#fff;cursor:default}.ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj{color:#eee;font-family:Roboto-light,arial,sans-serif;height:40px;line-height:40px}.ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS{background-color:#242223;float:left;font-family:Roboto-light,arial,sans-serif;font-size:12px;font-weight:500;padding-right:5px;text-transform:uppercase}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS{background-color:#323232;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;text-transform:none}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS{background:var(--dt-surface,#fff)}.ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf{margin-bottom:10px;padding-top:19px;width:100%}.ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe{border-top:1px solid #686868}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe{border-top:1px solid rgba(255,255,255,.15)}.ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc{color:#b6b6b6;font-size:12px;padding-bottom:20px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc{color:rgba(255,255,255,.57)}.ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b{display:inline-block;text-align:left;width:-moz-calc(100% - 150px);width:calc(100% - 150px)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b{color:rgba(255,255,255,.9);width:-moz-calc(100% - 128px);width:calc(100% - 128px)}.ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc{display:inline-block}.ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc.ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc{vertical-align:top;width:150px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc.ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc{width:128px}.ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc.ndfHFb-c4YZDc-MZArnb-BA389-V67aGc{width:-moz-calc(100% - 100px);width:calc(100% - 100px)}.ndfHFb-c4YZDc-MZArnb-P86uke-PntVL{display:inline-block;vertical-align:top;width:100%}.ndfHFb-c4YZDc-MZArnb-P86uke-Bz112c{float:left;margin-right:12px;margin-top:5px;width:16px;height:13px}.ndfHFb-c4YZDc-MZArnb-P86uke-hSRGPd{cursor:pointer;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.ndfHFb-c4YZDc-MZArnb-P86uke-hSRGPd:focus,.ndfHFb-c4YZDc-MZArnb-P86uke-hSRGPd:hover{text-decoration:underline}.ndfHFb-c4YZDc-MZArnb-BA389-V1ur5d{line-height:24px;margin-left:36px;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.ndfHFb-c4YZDc-MZArnb-BA389-nNAX0{display:inline-block;float:right;overflow-x:hidden}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-BA389-nNAX0{color:rgba(255,255,255,.9)}.ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c{line-height:24px;padding-bottom:10px}.ndfHFb-c4YZDc-MZArnb-Tswv1b-BKwaUc{-moz-box-sizing:content-box;box-sizing:content-box;border:none;width:100%}.ndfHFb-c4YZDc-MZArnb-ij8cu{font-weight:normal;padding-bottom:20px;word-wrap:break-word}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-ij8cu{margin-right:44px}.ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe{background-color:#242223;cursor:pointer;float:right;margin-top:8px;padding-left:3px}.ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:#242223;background-image:-moz-linear-gradient(top,#333,#222);background-image:linear-gradient(top,#333,#222)}.ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -760px;height:24px;width:24px}.ndfHFb-c4YZDc-MZArnb-ij8cu-DyVDA{-moz-box-sizing:border-box;box-sizing:border-box;min-height:75px;max-width:350px;overflow-y:auto;width:100%}.ndfHFb-c4YZDc-MZArnb-Tswv1b-nUpftc,.ndfHFb-c4YZDc-MZArnb-RDNXzf-nUpftc{-moz-user-select:text;padding:15px}.ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-bN97Pc-u0pjoe-fmcmS{font-size:12px;line-height:20px}.ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c{margin:1px 0}.ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c{float:left;height:24px}.ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c .ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c{height:24px;position:relative;width:24px}.ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e{background-color:#464445;-moz-border-radius:50%;border-radius:50%;display:inline-block;height:24px;width:24px}.ndfHFb-c4YZDc-MZArnb-ynfwJ-bF1uUb{color:#fff;line-height:24px;text-align:center;text-transform:uppercase;vertical-align:middle}.ndfHFb-c4YZDc-MZArnb-JNdkSc-YLEF4c{background-position:0 -2160px}.ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c{background-position:0 -2400px}.ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c-SfQLQb-hSRGPd{background-position:0 -280px}.ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c{background-position:0 -720px}.ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c-SfQLQb-hSRGPd{background-position:0 -480px}.ndfHFb-c4YZDc-MZArnb-YLEF4c-Bz112c{height:20px;margin:2px;width:20px}.ndfHFb-c4YZDc-MZArnb-nupQLb-BA389-Ne3sFf{display:inline-block}.ndfHFb-c4YZDc-MZArnb-MPu53c{-moz-box-sizing:border-box;box-sizing:border-box;border:2px solid #c1bfbf;-moz-border-radius:2px;border-radius:2px;cursor:pointer;float:right;height:20px;width:20px}.ndfHFb-c4YZDc-MZArnb-MPu53c-bN97Pc{height:16px}.ndfHFb-c4YZDc-MZArnb-MPu53c-fmcmS{font-size:20px;font-weight:bold;line-height:16px;position:absolute}.ndfHFb-c4YZDc-MZArnb-MPu53c-Bz112c{background-position:0 -1680px;display:inline-block;height:14px;width:14px;margin-top:2px;margin-left:1px}.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-MZArnb-b0t70b{width:100%;right:0;-moz-transition:right .218s cubic-bezier(0,0,0.2,1);transition:right .218s cubic-bezier(0,0,0.2,1)}.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-MZArnb-b0t70b-L6cTce{display:block;right:-100%;-moz-transition:right .218 cubic-bezier(0.4,0,1,1);transition:right .218 cubic-bezier(0.4,0,1,1)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -288px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-J2xVie-Bz112c{background-position:0 -3674px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-JNdkSc-YLEF4c{background-position:0 -3138px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c{background-position:0 -1264px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-QIk5de-YLEF4c-SfQLQb-hSRGPd{background-position:0 -816px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c{background-position:0 -168px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-nE4Pff-YLEF4c-SfQLQb-hSRGPd{background-position:0 -736px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe:not(.ndfHFb-c4YZDc-LgbsSe-ZmdkE){background-color:#323232;padding:8px;margin-top:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe:not(.ndfHFb-c4YZDc-LgbsSe-ZmdkE){background-color:transparent}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe{background-color:rgba(196,199,197,.12)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-TvD9Pc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{float:right;margin:8px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -3178px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-b0t70b .ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{margin-top:-8px}.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb{border-top:1px solid #686868;font-size:12px;font-weight:normal;outline:none;padding:18px 0 7px 0;position:relative;zoom:1}.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb:first-child{border-top-color:transparent}.ndfHFb-c4YZDc-MZArnb-jNm5if-haAclf{margin-left:55px}.ndfHFb-c4YZDc-MZArnb-jNm5if{min-height:48px;position:relative}.ndfHFb-c4YZDc-MZArnb-jNm5if-tJHJj{color:#757272;font-style:italic}.ndfHFb-c4YZDc-MZArnb-jNm5if-EieU8{background-color:#211f20;margin:4px 0 3px}.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb{margin-bottom:10px}.ndfHFb-c4YZDc-MZArnb-jNm5if-gqY2Od{color:#b6b6b6;display:inline-block;font-weight:bold;max-width:180px;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.ndfHFb-c4YZDc-MZArnb-jNm5if-IIEkAe .ndfHFb-c4YZDc-MZArnb-jNm5if-gqY2Od{max-width:120px}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-bN97Pc .ndfHFb-c4YZDc-MZArnb-jNm5if-gqY2Od{font-style:normal;margin-right:4px}.ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c{-moz-border-radius:50%;border-radius:50%;height:48px;left:0;position:absolute;width:48px}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb .ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c{-moz-border-radius:0;border-radius:0;height:24px;left:6px;width:24px}.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e{height:48px;width:48px;left:0;position:absolute}.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-ynfwJ-bF1uUb{font-size:24px;line-height:48px}.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb .ndfHFb-c4YZDc-MZArnb-zTETae-YLEF4c-JUCs7e{-moz-border-radius:0;border-radius:0;height:24px;width:24px}.ndfHFb-c4YZDc-MZArnb-jNm5if-pXBrqb .ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb .ndfHFb-c4YZDc-MZArnb-ynfwJ-bF1uUb{font-size:12px;line-height:24px}.ndfHFb-c4YZDc-MZArnb-jNm5if-biJjHb-haAclf{color:#c1bfbf;font-size:10px;padding-top:2px;position:absolute;right:0;top:0}.ndfHFb-c4YZDc-MZArnb-jNm5if-biJjHb{display:inline-block;padding:0 3px}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-bN97Pc .ndfHFb-c4YZDc-MZArnb-jNm5if-biJjHb{color:#c1bfbf;font-size:10px;padding:3px 0;position:relative}.ndfHFb-c4YZDc-MZArnb-jNm5if-bN97Pc{color:#fff;margin-top:5px;word-wrap:break-word;top:-7px;zoom:1}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb{border-top:1px solid #242223;color:#888;min-height:24px;padding:6px 3px 0 6px;position:relative}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb:first-child{border-top-color:transparent}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-bN97Pc{padding-left:30px}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-fmcmS{line-height:140%;position:relative;top:-3px;width:100%}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-qJTHM{color:#fff;display:inline;margin:0;position:relative;top:-4px;width:100%;word-wrap:break-word}.ndfHFb-c4YZDc-MZArnb-IIEkAe-jNm5if-Ne3sFf{display:inline;padding-right:18px}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-JIbuQc{color:#fff;display:inline;font-style:italic;position:relative;top:-4px}.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-JIbuQc+.ndfHFb-c4YZDc-MZArnb-jNm5if-xtcdFb-qJTHM{display:block}.ndfHFb-c4YZDc-MZArnb-IIEkAe-jNm5if-Bz112c{background-position:0 -1680px;display:inline-block;height:12px;margin-left:3px;position:absolute;right:0;width:15px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-IIEkAe-jNm5if-Bz112c{background-position:0 -2504px}.ndfHFb-c4YZDc-C7uZwb-LgbsSe .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{filter:alpha(opacity=87);opacity:0.87;margin-left:auto;margin-right:auto;margin-top:3px;height:21px;width:21px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{filter:alpha(opacity=87);opacity:0.87;margin-right:auto;margin-top:3px;height:21px;width:21px}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-C7uZwb-LgbsSe-SfQLQb-Bz112c.ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{filter:alpha(opacity=47);opacity:0.47}.ndfHFb-c4YZDc-C7uZwb-LgbsSe-SfQLQb-Bz112c.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-nupQLb-Bz112c{background-position:0 -1040px}.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c{background-position:0 -1880px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c{background-position:0 -1560px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-nupQLb-Bz112c{background-position:0 -2480px}.ndfHFb-c4YZDc-VkLyEc-Bz112c{background-position:0 -2320px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-VkLyEc-Bz112c{background-position:0 -1480px}.ndfHFb-c4YZDc-euCgFf-Bz112c{background-position:0 -1440px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-euCgFf-Bz112c{background-position:0 -1200px}.ndfHFb-c4YZDc-hN7jy-Bz112c{background-position:0 -2200px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-hN7jy-Bz112c{background-position:0 -2280px}.ndfHFb-c4YZDc-PEFSMe-Bz112c{background-position:0 -2240px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-PEFSMe-Bz112c{background-position:0 -360px}.ndfHFb-c4YZDc-uQPRwe-uWtm3-Bz112c{background-position:0 -1800px}.ndfHFb-c4YZDc-w37qKe-Bz112c{background-position:0 -440px}.ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c{background-position:0 -40px}.ndfHFb-c4YZDc-Vkfede-fI6EEc-Bz112c{background-position:0 -1720px}.ndfHFb-c4YZDc-J2Tr8e-fI6EEc-Bz112c{background-position:0 -2000px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg');background-size:auto;margin-left:2px;left:8px;top:3px}.ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{top:2px}.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c.ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c,.ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c.ndfHFb-c4YZDc-w37qKe-Bz112c{height:24px;margin-left:0;margin-top:-1px;width:24px}.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe{border:1px solid #1a73e8;-moz-border-radius:2px;border-radius:2px;-moz-box-shadow:inset 0 1px 0 rgba(101,101,101,.1);box-shadow:inset 0 1px 0 rgba(101,101,101,.1);background-color:#1a73e8;color:#fff;display:inline-block;font-size:11px;font-weight:bold;text-align:center;text-shadow:0 1px 0 rgba(0,0,0,.8);height:28px;line-height:28px;margin-top:20px;min-width:54px;padding:0 20px 0 7px;vertical-align:middle;white-space:nowrap}.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg');height:21px;margin-top:4px;position:absolute;width:21px}.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-fmcmS{margin-left:35px;margin-right:10px}.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe{background-color:#1a73e8;background-image:-moz-linear-gradient(top,#1a73e8,#357ae8);background-image:linear-gradient(top,#1a73e8,#357ae8)}.ndfHFb-c4YZDc-LgbsSe-auswjd.ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe{-moz-box-shadow:inset 0 1px 6px rgba(0,0,0,.8);box-shadow:inset 0 1px 6px rgba(0,0,0,.8)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-C7uZwb-LgbsSe .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{margin-top:0;height:24px;width:24px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{margin-top:0;height:24px;width:24px;background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg')}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-bN97Pc-nupQLb-LgbsSe-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg')}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nupQLb-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nupQLb-Bz112c{background-position:0 -2384px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c{background-position:0 -408px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c{background-position:0 -3530px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-FNFY6c-bEDTcc-oxvKad-Bz112c{background-position:0 -408px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-nupQLb-Bz112c{background-position:0 -2384px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-nupQLb-Bz112c{background-position:0 -632px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-VkLyEc-Bz112c{background-position:0 -2584px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-VkLyEc-Bz112c{background-position:0 -2890px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-VkLyEc-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-VkLyEc-Bz112c{background-position:0 -2584px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-euCgFf-Bz112c{background-position:0 -3218px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-euCgFf-Bz112c{background-position:0 -2994px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-euCgFf-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-euCgFf-Bz112c{background-position:0 -3218px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-hN7jy-Bz112c{background-position:0 -2016px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-hN7jy-Bz112c{background-position:0 -1368px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-hN7jy-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-hN7jy-Bz112c{background-position:0 -2016px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c{background-position:0 -3258px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c{background-position:0 -1856px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-dMDEpe-tgaKEf-Bz112c{background-position:0 -3258px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-PEFSMe-Bz112c{background-position:0 -3426px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-PEFSMe-Bz112c{background-position:0 -512px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-PEFSMe-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-PEFSMe-Bz112c{background-position:0 -3426px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-uQPRwe-uWtm3-Bz112c{background-position:0 -3098px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-uQPRwe-uWtm3-Bz112c{background-position:0 -3714px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-w37qKe-Bz112c{background-position:0 -1200px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-w37qKe-Bz112c{background-position:0 -1568px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c{background-position:0 -672px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-ndfHFb-w37qKe-Bz112c{background-position:0 -328px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Vkfede-fI6EEc-Bz112c{background-position:0 -2930px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Vkfede-fI6EEc-Bz112c{background-position:0 -1672px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-J2Tr8e-fI6EEc-Bz112c{background-position:0 -88px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-J2Tr8e-fI6EEc-Bz112c{background-position:0 -1488px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-Bz112c{background-position:0 -1712px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-Bz112c{background-position:0 -208px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-GSQQnc-LgbsSe{background-position:0 -368px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-GSQQnc-LgbsSe{background-position:0 -2304px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c{background-position:0 -2602px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3338px;transform:scale(0.8) translateX(3px) translateY(9px);width:24px;height:24px;pointer-events:none}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-hOcTPc .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c{transform:scale(0.8);margin-left:4px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-RDNXzf-OWB6Me-Bz112c{background-position:0 -40px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c{background-position:0 -1632px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-htvI8d-jNm5if-Bz112c{background-position:0 -2602px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-ge6pde-Bz112c .ndfHFb-aZ2wEe{display:block}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-pGuBYc-Bz112c{background-position:0 -472px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-MqcBrc-Bz112c{background-position:0 -3634px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-MqcBrc-Bz112c{background-position:0 -2850px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-SjW3R-Bz112c{background-position:0 -3034px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-SjW3R-Bz112c{background-position:0 -2970px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-lCdvJf-Bz112c{background-position:0 -1896px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c.ndfHFb-c4YZDc-lCdvJf-Bz112c{background-position:0 -128px}.ndfHFb-c4YZDc-E90Ek{background-color:rgba(0,0,0,.75);display:inline-block;margin-right:50px;padding:2px;width:500px}.ndfHFb-c4YZDc-E90Ek-tJHJj{font-size:18px;margin:10px;text-align:center}.ndfHFb-c4YZDc-E90Ek-LgbsSe{background-color:dimgray;cursor:pointer;float:right;padding:10px}.ndfHFb-c4YZDc-E90Ek-bN97Pc{max-height:600px;max-width:600px;overflow-x:scroll}.ndfHFb-c4YZDc-E90Ek-Tswv1b-tJHJj{margin:10px;text-align:left}.ndfHFb-c4YZDc-E90Ek-Tswv1b-lTBxed{color:white;margin:0 10px}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe,.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center;position:absolute;z-index:2;pointer-events:all}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-B8qYne,.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-B8qYne,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-B8qYne{height:100%;width:100%;display:none;align-items:center;position:absolute;z-index:2;pointer-events:all}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-B8qYne-RJLb9c,.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-B8qYne-RJLb9c,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-B8qYne-RJLb9c{max-width:100%;max-height:100%}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-WbpZL,.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-WbpZL,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-WbpZL{height:100%;width:100%;display:none;align-items:center;z-index:2;pointer-events:all;background:#e8f0fe;color:#185abc;border:1px solid #185abc;-moz-border-radius:4px;border-radius:4px;box-sizing:border-box;cursor:pointer}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-jf2N7b-dIxMhd-zUk4Qd,.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-jf2N7b-dIxMhd-zUk4Qd,.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-jf2N7b-dIxMhd-zUk4Qd,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-jf2N7b-dIxMhd-zUk4Qd{height:100%;width:100%;display:none;align-items:center;z-index:2;pointer-events:all;background:#f1f3f4;color:#c0c0c0;border:1px solid #c0c0c0;-moz-border-radius:4px;border-radius:4px;box-sizing:border-box}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-jf2N7b-dIxMhd-MFS4be,.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-jf2N7b-dIxMhd-MFS4be,.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-jf2N7b-dIxMhd-MFS4be,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-jf2N7b-dIxMhd-MFS4be{height:100%;width:100%;display:none;align-items:center;z-index:2;pointer-events:all;background:transparent;color:#c0c0c0;border:1px solid #c0c0c0;-moz-border-radius:4px;border-radius:4px;box-sizing:border-box}.ndfHFb-c4YZDc-dZssN-yrriRe-JbbQac-LgbsSe{position:absolute;right:0;top:0;background:#3c4043;opacity:.4;-moz-border-radius:50%;border-radius:50%;display:none;height:24px;width:24px;pointer-events:all;z-index:2;cursor:pointer}.ndfHFb-c4YZDc-dZssN-yrriRe-JbbQac-LgbsSe-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3362px;height:11.62px;width:11.67px;margin:auto}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-WbpZL-fmcmS,.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-WbpZL-fmcmS,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-WbpZL-fmcmS{color:#174ea6;font-family:"Roboto Mono",monospace;font-style:normal;font-weight:bold;font-size:16px;line-height:22px;position:absolute;top:auto;bottom:auto;left:9.41%;right:78%}.ndfHFb-c4YZDc-dZssN-mKZypf-qFWjAd-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -2786px;height:13.33px;width:13.29px;position:absolute;top:auto;bottom:auto;right:14.31%}.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;align-items:center;position:absolute;z-index:2;pointer-events:all}.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-fmcmS{display:none;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:22px;line-height:20px;color:black}.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-suEOdc{position:absolute;background-color:#202124;color:#dadce0;font-family:"Roboto";font-style:normal;font-weight:400;font-size:14px;line-height:20px;letter-spacing:.2px;-moz-border-radius:4px;border-radius:4px;visibility:hidden;width:210px;height:max-content;top:42px;left:20px;padding:9px 13px}.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe:hover .ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-suEOdc{position:absolute;visibility:visible}.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe:hover{z-index:100}.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-FVVVue-WAutxc-zUk4Qd{display:none;width:100%;height:100%;align-items:center;background-color:#e8f0fe;color:#174ea6;position:absolute;z-index:2;pointer-events:all}.ndfHFb-c4YZDc-dZssN-B8qYne-gElRsf-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -2136px;height:17.61px;width:16px;position:absolute;top:auto;bottom:auto;left:18.5px;transform:scale(0.9375,0.9432)}.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-FVVVue-WAutxc-zUk4Qd,.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-FVVVue-WAutxc-zUk4Qd,.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-FVVVue-WAutxc-zUk4Qd{display:none;width:100%;height:100%;align-items:center;background-color:#e8f0fe;color:#174ea6;position:absolute;z-index:2;pointer-events:all}.ndfHFb-c4YZDc-dZssN-ikE8I-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -1608px;height:17.61px;width:16px;position:absolute;top:auto;bottom:auto;left:18.5px;transform:scale(0.9375,0.9432)}.ndfHFb-c4YZDc-dZssN-Wqqruc-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3506px;height:24px;width:24px;position:absolute;top:auto;bottom:auto;left:18.5px;transform:scale(0.9375,0.9432)}.ndfHFb-c4YZDc-dZssN-tekGAe-V1ur5d-yrriRe-FVVVue-WAutxc-zUk4Qd-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -1792px;height:17.61px;width:16px;position:absolute;top:auto;bottom:auto;left:18.5px;transform:scale(0.9375,0.9432)}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:0;outline:none;position:absolute;width:453px;background:#fff;-moz-box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);-moz-border-radius:8px;border-radius:8px;z-index:1194}.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:0;outline:none;position:absolute;width:340px;background:#fff;-moz-box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);-moz-border-radius:8px;border-radius:8px;z-index:1194}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:0;outline:none;position:absolute;width:468px;background:#fff;-moz-box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);-moz-border-radius:8px;border-radius:8px;z-index:1194}.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:0;outline:none;position:absolute;width:300px;background:#fff;-moz-box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);-moz-border-radius:8px;border-radius:8px;z-index:1194}.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:0;outline:none;position:absolute;width:350px;background:#fff;-moz-box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);-moz-border-radius:8px;border-radius:8px;z-index:1194}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-xJ5Hnf,.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-xJ5Hnf,.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-xJ5Hnf,.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-xJ5Hnf,.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-xJ5Hnf{background-color:#000;height:100%;left:0;position:fixed;top:0;width:100%;z-index:1194}.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe-xJ5Hnf{background-color:#000;height:100%;left:0;position:fixed;top:0;width:100%;z-index:1194}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-r4nke{margin:0 auto}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-r4nke,.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-r4nke,.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-r4nke,.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-r4nke{margin:24px 24px}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-r4nke-fmcmS,.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-r4nke-fmcmS,.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-r4nke-fmcmS,.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-r4nke-fmcmS,.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-r4nke-fmcmS{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;letter-spacing:0;line-height:1.75rem;color:#202124}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-HiaYvf{width:125px;height:125px;margin-bottom:33px;margin-top:39px;margin-right:auto;margin-left:auto;display:block}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-bN97Pc{letter-spacing:.01428571em;font-family:Roboto,Arial,sans-serif;font-size:.875rem;font-weight:400;line-height:1.25rem;color:#5f6368;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;justify-content:space-between;margin:16px 24px 12px;text-align:center}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-bN97Pc{color:#5f6368;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;justify-content:space-between;margin:0 12px 12px;text-align:left}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-g7W7Ed{color:#5f6368;font-family:"Roboto";font-style:normal;font-weight:400;font-size:14px;line-height:20px;letter-spacing:.2px;margin-bottom:22.6px;width:428px}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-MPu53c-bN97Pc{color:#3c4043;font-family:"Roboto";font-style:normal;font-weight:700;font-size:14px;line-height:20px;letter-spacing:.2px;text-align:left}.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-bN97Pc{letter-spacing:.01428571em;font-family:Roboto,Arial,sans-serif;font-size:.875rem;font-weight:400;line-height:1.25rem;color:#5f6368;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;justify-content:space-between;margin:16px 24px 12px;text-align:center}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-bN97Pc-PLDbbf{text-decoration:none;color:#1a73e8}.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-bN97Pc{letter-spacing:.01428571em;font-family:Roboto,Arial,sans-serif;font-size:.875rem;font-weight:400;line-height:1.25rem;color:#5f6368;justify-content:space-between;margin-top:0;margin-left:24px;margin-right:24px;margin-bottom:0;max-width:300px;overflow-wrap:break-word;text-align:center}.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-bN97Pc{color:#5f6368;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;justify-content:space-between;text-align:center}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-LgbsSe,.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-LgbsSe,.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-IbE0S-LgbsSe,.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-IbE0S-LgbsSe,.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-LgbsSe{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;line-height:20px;background:#fff;border:1px solid #dadce0;-moz-border-radius:4px;border-radius:4px;box-sizing:border-box;color:#1a73e8;margin:0 12px;min-width:70px;outline:none;padding:8px 24px;text-align:center;cursor:pointer}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-Wh8OAb-LgbsSe{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;line-height:20px;border:none;background:#1a73e8;box-sizing:border-box;-moz-border-radius:4px;border-radius:4px;color:#fff;margin:0 12px;min-width:70px;outline:none;padding:8px 24px;text-align:center;cursor:pointer;opacity:30%}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-Wh8OAb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-qnnXGd{opacity:100%}.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-ERydpb-LgbsSe{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;line-height:20px;border:none;background:#d93025;box-sizing:border-box;-moz-border-radius:4px;border-radius:4px;color:#fff;margin:0 12px;min-width:70px;outline:none;padding:8px 24px;text-align:center;cursor:pointer}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-HiaYvf{width:97px;height:97px;margin-bottom:36px;margin-right:auto;margin-left:auto}.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-c6xFrd{margin:21px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;padding:0}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-c6xFrd,.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-c6xFrd{margin-left:auto;margin-right:auto;margin-bottom:18px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row}.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-c6xFrd{margin-right:22px;margin-left:auto;margin-bottom:18px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;padding:0}.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-c6xFrd{margin-top:22px;margin-right:22px;margin-left:auto;margin-bottom:18px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;padding:0}.ndfHFb-c4YZDc-dZssN-udLbKb-Sx9Kwc-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-Wh8OAb-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-Dogjgd-eKpHRd-UDALgf-Sx9Kwc-IbE0S-LgbsSe .ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-u0pjoe-Sx9Kwc-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-ERydpb-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-ERydpb-eizL8e-Sx9Kwc-IbE0S-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-ERydpb-udLbKb-Sx9Kwc-LgbsSe:hover{cursor:pointer}.ndfHFb-c4YZDc-dZssN-ORHb-haAclf{position:relative;top:0;z-index:3}.ndfHFb-c4YZDc-dZssN-ORHb-r4nke{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.125rem;font-weight:400;letter-spacing:0;line-height:1.5rem;-moz-border-radius:0;border-radius:0;background-color:#000;color:#fff;padding-left:24px;height:56px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-r4nke{height:64px}.ndfHFb-c4YZDc-dZssN-ORHb{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;letter-spacing:.00625em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1rem;font-weight:500;line-height:1.5rem;background-color:#e8f0fe;-moz-border-radius:0;border-radius:0;color:#202124;height:48px;width:100%;-moz-box-shadow:0px 1px 2px 0px rgba(60,64,67,.30),0px 2px 6px 2px rgba(60,64,67,.15);box-shadow:0px 1px 2px 0px rgba(60,64,67,.30),0px 2px 6px 2px rgba(60,64,67,.15)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb{background:#7cacf8}.ndfHFb-c4YZDc-dZssN-ORHb-bN97Pc{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;justify-content:space-between;width:100%}.ndfHFb-c4YZDc-dZssN-ORHb-Ne3sFf{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-Ne3sFf{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-dZssN-ORHb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -712px;height:16px;margin:0 13px 0 25px;width:18px;transform:scale(1.076,1)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-Bz112c{background-position:0 -976px;height:24px;margin:0 16px;width:24px}.ndfHFb-c4YZDc-dZssN-ORHb-LQLjdd{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-flex:none;flex:none;box-flex:0;flex-grow:0;margin:8px 0;-moz-box-ordinal-group:0;order:0}.ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe,.ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe{color:#1a73e8;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;-moz-border-radius:5px;border-radius:5px;letter-spacing:.25px;line-height:20px;text-align:center;text-decoration:none;margin:0 12px;padding:6px 14px;cursor:pointer}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe{color:#202124;background:transparent;font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em)}.ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe:hover{background:#f8fbff}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-LgbsSe:hover,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-LgbsSe:hover,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe:hover{background:transparent}.ndfHFb-c4YZDc-dZssN-ORHb-LgbsSe-L6cTce{display:none}.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe{color:#fff;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;-moz-border-radius:5px;border-radius:5px;letter-spacing:.25px;line-height:20px;text-align:center;text-decoration:none;margin:0 12px;padding:6px 14px;background-color:#1a73e8;cursor:pointer;opacity:30%;pointer-events:none}.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe:hover{background:#2b7de9}.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-sM5MNb,.ndfHFb-c4YZDc-dZssN-ORHb-ERydpb-sM5MNb,.ndfHFb-c4YZDc-dZssN-ORHb-nUpftc-MZArnb-sM5MNb{background:none}.ndfHFb-c4YZDc-dZssN-ORHb-SYOSDb-SDqDXe-LgbsSe.ndfHFb-c4YZDc-LgbsSe-qnnXGd{opacity:100%;pointer-events:auto}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-haAclf{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;letter-spacing:.00625em;font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1rem;font-weight:500;line-height:1.5rem;background-color:#e8f0fe;-moz-border-radius:0;border-radius:0;color:#202124;height:48px;width:100%;-moz-box-shadow:0px 1px 2px 0px rgba(60,64,67,.30),0px 2px 6px 2px rgba(60,64,67,.15);box-shadow:0px 1px 2px 0px rgba(60,64,67,.30),0px 2px 6px 2px rgba(60,64,67,.15)}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-bN97Pc{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;justify-content:space-between;width:100%}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Ne3sFf{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -712px;height:16px;margin:0 13px 0 25px;width:18px;transform:scale(1.076,1)}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-LQLjdd{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-box-flex:none;flex:none;box-flex:0;flex-grow:0;margin:8px 0;-moz-box-ordinal-group:0;order:0}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-LgbsSe,.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-LgbsSe{color:#1a73e8;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;-moz-border-radius:5px;border-radius:5px;letter-spacing:.25px;line-height:20px;text-align:center;text-decoration:none;margin:0 12px;padding:6px 14px;cursor:pointer}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-LgbsSe:hover,.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-LgbsSe:hover{background:#f8fbff}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-LgbsSe{color:#fff;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;-moz-border-radius:5px;border-radius:5px;letter-spacing:.25px;line-height:20px;text-align:center;text-decoration:none;margin:0 12px;padding:6px 14px;background-color:#1a73e8;cursor:pointer}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-LgbsSe:hover{background:#2b7de9}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-mKZypf-sM5MNb,.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-ERydpb-sM5MNb,.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-nUpftc-MZArnb-sM5MNb{background:none}.ndfHFb-c4YZDc-dZssN-FVVVue-ORHb-haAclf.ndfHFb-c4YZDc-ORHb-L6cTce{display:none}.ndfHFb-c4YZDc-dZssN-x5yx9d-b0t70b{background:white;bottom:0;position:absolute;right:0;top:0;display:none}.ndfHFb-c4YZDc-dZssN-x5yx9d-L5Fo6c{border:none;height:100%;width:100%}.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe{width:100%;height:100%;top:50%}.ndfHFb-c4YZDc-EglORb-ge6pde.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe{min-width:0}.ndfHFb-c4YZDc-dZssN-ge6pde-aZ2wEe-haAclf{z-index:9000}.ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c{background-repeat:no-repeat;filter:alpha(opacity=87);opacity:0.87;margin-left:auto;margin-right:auto;margin-top:3px;height:21px;width:19px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-PlOyMe-bN97Pc{line-height:32px}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/v-spinner_dark.gif')}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me.ndfHFb-c4YZDc-Wrql6b-PlOyMe{background-color:transparent}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c:not([onclick]):not(:link):not(:visited){background-image:none;height:21px;width:21px}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c:not([onclick]):not(:link):not(:visited){background-image:none;height:24px;width:24px}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c .ndfHFb-aZ2wEe{display:block}.ndfHFb-c4YZDc-cnqxLd{background-color:#121212;bottom:0;color:#fff;font-size:0;height:0;position:absolute;-moz-transition:height .218s ease-out;transition:height .218s ease-out;width:100%;z-index:2}.ndfHFb-c4YZDc-cnqxLd-SmKAyb{overflow-x:auto;overflow-y:hidden;position:absolute;top:0;width:100%;white-space:nowrap}.ndfHFb-c4YZDc-cnqxLd-OEVmcd{border:3px solid #fff;-moz-border-radius:3px;border-radius:3px;position:absolute;height:63px;width:84px;margin-top:3px}.ndfHFb-c4YZDc-cnqxLd-LQLjdd{position:absolute;height:25px;z-index:1}.ndfHFb-c4YZDc-cnqxLd-LQLjdd-hOcTPc{left:12px}.ndfHFb-c4YZDc-cnqxLd-LQLjdd-AeOLfc{right:12px}.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe{background-color:rgba(0,0,0,.2);-moz-border-radius:3px;border-radius:3px;color:rgba(255,255,255,0.87);font-size:11px;text-align:center;text-shadow:0 1px 1px rgba(0,0,0,.8);height:25px;line-height:25px;padding:0 13px}.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:rgba(0,0,0,.4)}.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe-IwzHHe,.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-cnqxLd-N7Eqid-bF1uUb{background-color:rgba(0,0,0,.6)}.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE,.ndfHFb-c4YZDc-cnqxLd-LQLjdd .ndfHFb-c4YZDc-cnqxLd-N7Eqid-bF1uUb.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:rgba(0,0,0,.9)}.ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c{background-position:0 -1080px;display:inline-block;height:21px;margin-right:4px;vertical-align:top;width:21px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c{background-position:0 -2160px}.ndfHFb-c4YZDc-cnqxLd-LSZ0mb.ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c{background-position:0 -960px;height:16px;margin-top:5px;padding-left:5px;width:16px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-cnqxLd-LSZ0mb.ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-cnqxLd-LSZ0mb-Bz112c{background-position:0 -1936px}.ndfHFb-c4YZDc-cnqxLd-LSZ0mb-fmcmS{display:inline-block;margin-top:1px;vertical-align:middle}.ndfHFb-c4YZDc-n5VRYe-ma6Yeb,.ndfHFb-c4YZDc-n5VRYe-AeOLfc,.ndfHFb-c4YZDc-n5VRYe-cGMI2b,.ndfHFb-c4YZDc-n5VRYe-hOcTPc{z-index:1;position:absolute}.ndfHFb-c4YZDc-n5VRYe-ma6Yeb,.ndfHFb-c4YZDc-n5VRYe-cGMI2b{height:8px;left:0;right:0}.ndfHFb-c4YZDc-n5VRYe-AeOLfc,.ndfHFb-c4YZDc-n5VRYe-hOcTPc{bottom:0;top:0;width:8px}.ndfHFb-c4YZDc-n5VRYe-ma6Yeb{background-color:none;background-image:-moz-linear-gradient(top,rgba(0,0,0,.35),rgba(0,0,0,0));background-image:linear-gradient(top,rgba(0,0,0,.35),rgba(0,0,0,0));top:0}.ndfHFb-c4YZDc-n5VRYe-AeOLfc{background-color:none;background-image:-moz-linear-gradient(right,rgba(0,0,0,.35),rgba(0,0,0,0));background-image:linear-gradient(right,rgba(0,0,0,.35),rgba(0,0,0,0));right:0}.ndfHFb-c4YZDc-n5VRYe-cGMI2b{background-color:none;background-image:-moz-linear-gradient(bottom,rgba(0,0,0,.35),rgba(0,0,0,0));background-image:linear-gradient(bottom,rgba(0,0,0,.35),rgba(0,0,0,0));bottom:0}.ndfHFb-c4YZDc-n5VRYe-hOcTPc{background-color:none;background-image:-moz-linear-gradient(left,rgba(0,0,0,.35),rgba(0,0,0,0));background-image:linear-gradient(left,rgba(0,0,0,.35),rgba(0,0,0,0));left:0}.ndfHFb-c4YZDc-Sx9Kwc.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc{padding:0}.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde{background-color:#f3f3f3;height:100%;position:relative;width:100%}.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde .ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-Sx9Kwc-ge6pde-k4Qmrd{text-align:center;width:100%;position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-t2cHAd-DWWcKd-ZpdDCc-ge6pde-RJLb9c{background-image:url('//ssl.gstatic.com/ui/v1/activityindicator/loading_bg_f5.gif');background-repeat:no-repeat;display:inline-block;height:19px;position:relative;top:3px;width:19px}.ndfHFb-c4YZDc-w5vlXd{border:1px solid transparent}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg')!important;background-repeat:no-repeat}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg')!important}.ndfHFb-c4YZDc-L5Fo6c-nUpftc{position:absolute}.ndfHFb-c4YZDc-HiaYvf{position:absolute;background-color:white;background-image:-moz-linear-gradient(45deg,#efefef 25%,transparent 25%,transparent 75%,#efefef 75%,#efefef),-moz-linear-gradient(45deg,#efefef 25%,transparent 25%,transparent 75%,#efefef 75%,#efefef);background-image:linear-gradient(45deg,#efefef 25%,transparent 25%,transparent 75%,#efefef 75%,#efefef),linear-gradient(45deg,#efefef 25%,transparent 25%,transparent 75%,#efefef 75%,#efefef);background-position:0 0,10px 10px;-moz-background-size:21px 21px;background-size:21px 21px;-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);-moz-user-select:none}.ndfHFb-c4YZDc-HiaYvf-s2gQvd{bottom:0;left:0;overflow:auto;position:absolute;right:0;top:0}.ndfHFb-c4YZDc-HiaYvf-s2gQvd .ndfHFb-c4YZDc-wvGCSb-gkA7Yd{right:initial}.ndfHFb-c4YZDc-HiaYvf-haAclf .ndfHFb-c4YZDc-TvD9Pc-qnnXGd,.ndfHFb-c4YZDc-HiaYvf-RJLb9c{height:100%;position:absolute;width:100%}.ndfHFb-c4YZDc-HiaYvf.ndfHFb-c4YZDc-HiaYvf-gvZm2b-qnnXGd{cursor:crosshair}.ndfHFb-c4YZDc-HiaYvf-lI7fHe-oYxtQd{-moz-box-shadow:0px 2px 4px 0px rgba(0,0,0,.5);box-shadow:0px 2px 4px 0px rgba(0,0,0,.5);-moz-border-radius:3px;border-radius:3px;position:absolute;z-index:1}.ndfHFb-c4YZDc-HiaYvf-gvZm2b{-moz-box-shadow:0px 2px 4px 0px rgba(0,0,0,.5);box-shadow:0px 2px 4px 0px rgba(0,0,0,.5);-moz-border-radius:3px;border-radius:3px;position:absolute}.ndfHFb-c4YZDc-HiaYvf-AHUcCb-oYxtQd.ndfHFb-c4YZDc-HiaYvf-lI7fHe-oYxtQd,.ndfHFb-c4YZDc-HiaYvf-gvZm2b{z-index:2}.ndfHFb-c4YZDc-HiaYvf-gvZm2b-SmKAyb,.ndfHFb-c4YZDc-HiaYvf-gvZm2b-n0tgWb{left:0;top:0;right:0;bottom:0;position:absolute}.ndfHFb-c4YZDc-HiaYvf-gvZm2b-SmKAyb{-moz-border-radius:2px;border-radius:2px;border:2px solid #fff;margin:1px;z-index:1}.ndfHFb-c4YZDc-HiaYvf-gvZm2b-n0tgWb{-moz-border-radius:3px;border-radius:3px;border:2px solid rgba(243,179,0,.5);z-index:2}.ndfHFb-c4YZDc-HiaYvf-mvZqyf{width:100%;height:100%;position:absolute;border:30000px solid #000;-moz-border-radius:30003px;border-radius:30003px;transform:translate(-30000px,-30000px);opacity:0;transition:opacity .4s ease;pointer-events:none}.ndfHFb-c4YZDc-HiaYvf-AHUcCb-oYxtQd .ndfHFb-c4YZDc-HiaYvf-mvZqyf,.ndfHFb-c4YZDc-HiaYvf-gvZm2b .ndfHFb-c4YZDc-HiaYvf-mvZqyf{opacity:.5}.ndfHFb-c4YZDc-RDNXzf-L6cTce .ndfHFb-c4YZDc-HiaYvf-lI7fHe-oYxtQd{display:none}.ndfHFb-c4YZDc-dkyuHd-ostUZ{position:absolute;min-width:400px;max-width:568px;line-height:20px;top:8px;background:#1a73e8;color:white;overflow:hidden;-moz-border-radius:2px;border-radius:2px;transform:translate(-50%,-64px);display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;align-items:center;-moz-box-shadow:0px 2px 4px rgba(0,0,0,.5);box-shadow:0px 2px 4px rgba(0,0,0,.5);-moz-transition:transform 0.15s;transition:transform 0.15s;z-index:4;left:50%}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ{background:#7cacf8;-moz-border-radius:8px;border-radius:8px;min-width:364px;-moz-box-shadow:none;box-shadow:none;color:#000;font:var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-title-medium-spacing,0.00625em);justify-content:space-between}.ndfHFb-c4YZDc-dkyuHd-ostUZ.ndfHFb-c4YZDc-dkyuHd-ostUZ-TSZdd{height:auto;transform:translate(-50%,0px)}.ndfHFb-c4YZDc-dkyuHd-ostUZ-Ne3sFf{padding:10px 32px 10px 16px;font-size:14px;font-weight:500;float:left}.ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S,.ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:visited{margin-left:auto;margin-top:auto;margin-bottom:auto;text-transform:uppercase;font-size:14px;cursor:pointer;padding:10px 16px;text-decoration:none;float:right}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:visited{text-transform:none;width:24px;height:24px}.ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S.ndfHFb-c4YZDc-LgbsSe-XpnDCe,.ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:hover{outline:white auto 5px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S .ndfHFb-c4YZDc-Bz112c{background-position:0 -3570px;width:24px;height:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S.ndfHFb-c4YZDc-LgbsSe-XpnDCe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-dkyuHd-ostUZ-IbE0S:hover{outline:none}.ndfHFb-c4YZDc-oKVyEf-haAclf,.ndfHFb-c4YZDc-oKVyEf-haAclf .ndfHFb-c4YZDc-TvD9Pc-qnnXGd{height:100%;position:absolute;width:100%}.ndfHFb-c4YZDc-oKVyEf-s2gQvd{bottom:0;left:0;overflow:auto;position:absolute;right:0;top:0}.ndfHFb-c4YZDc-oKVyEf-s2gQvd .ndfHFb-c4YZDc-wvGCSb-gkA7Yd{right:initial}@media print{.ndfHFb-c4YZDc-oKVyEf-PEFSMe-OWB6Me{display:none}}.ndfHFb-c4YZDc-LzGo7c{display:inline-block;font-size:12px;margin-bottom:10px;margin-left:5px;opacity:.7}.ndfHFb-c4YZDc-LzGo7c-fmcmS{color:#fff;display:inline-block;margin-right:4px}.ndfHFb-c4YZDc-hSRGPd-LgbsSe{color:#b3b3b3;cursor:pointer;text-decoration:underline}.ndfHFb-c4YZDc-xl07Ob,.ndfHFb-c4YZDc-mg9Pef{-moz-box-shadow:0 2px 4px rgba(0,0,0,.2);box-shadow:0 2px 4px rgba(0,0,0,.2);background:#fff;color:#333;font-family:arial,sans-serif;font-size:13px;border:1px solid #919191;line-height:18px;overflow-y:auto;position:absolute;z-index:1293;outline:1px solid transparent}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-xl07Ob,.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-mg9Pef{-moz-box-shadow:0 4px 8px rgba(0,0,0,.35);box-shadow:0 4px 8px rgba(0,0,0,.35);font-family:"Google Sans",Roboto,arial,sans-serif;border:0;-moz-border-radius:2px;border-radius:2px;line-height:34px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-xl07Ob,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-mg9Pef{background:var(--dt-surface,#fff);-moz-border-radius:4px;border-radius:4px}.ndfHFb-c4YZDc-j7LFlb{cursor:pointer;list-style:none;padding:6px 6em 6px 37px;position:relative;white-space:nowrap}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb{padding:1px 60px 1px 52px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb{padding-top:0;padding-bottom:0;height:34px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center}.ndfHFb-c4YZDc-j7LFlb-Bz112c{background-size:contain;height:16px;left:10px;position:absolute;top:6px;width:16px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-Bz112c{left:16px;height:20px;width:20px}.ndfHFb-c4YZDc-j7LFlb-sn54Q{background-color:#f1f1f1;border-color:#f1f1f1;border-style:dotted;border-width:1px 0;padding:5px 6em 5px 37px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-sn54Q{background-color:#dfdfdf;border-color:#dfdfdf;padding:0 60px 0 52px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb-sn54Q{background:#373737;border:none}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb:hover{background:#2f2f2f;border:none}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb:focus,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-j7LFlb:active{background:#373737;border:none}.ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c{top:5px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c{top:6px}.ndfHFb-c4YZDc-xl07Ob-tJHJj{color:#595959;cursor:default;font-size:12px;list-style:none;padding:6px 6em 6px 6px;position:relative;white-space:nowrap}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-tJHJj{padding:0 24px 0 12px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-tJHJj{color:var(--dt-on-surface,#3c4043)}.ndfHFb-c4YZDc-xl07Ob-hgDUwe{border-bottom:1px solid #444}.ndfHFb-c4YZDc-xl07Ob-WfNeFe-tJHJj{background-color:#efefef;font-style:italic}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-hgDUwe{border-color:#dfdfdf;margin:8px 0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-xl07Ob-hgDUwe{border-color:var(--dt-outline-variant,#dadce0);margin:8px 0}.ndfHFb-c4YZDc-mg9Pef .ndfHFb-c4YZDc-j7LFlb{line-height:36px;padding:0 40px 0 16px}.ndfHFb-c4YZDc-mg9Pef .ndfHFb-c4YZDc-j7LFlb-sn54Q{border:none;color:rgba(0,0,0,.7)}.ndfHFb-c4YZDc-mg9Pef{padding:8px 0}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-j7LFlb-bN97Pc{color:var(--dt-on-surface,#3c4043);font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-j7LFlb-bN97Pc .ndfHFb-c4YZDc-Bz112c{transform:scale(0.83)}.ndfHFb-c4YZDc-EglORb-haAclf{background-color:#4c494c;-moz-border-radius:12px;border-radius:12px;color:#fff;margin-bottom:40px;padding:20px;text-align:center;-moz-box-shadow:0px 10px 12px 5px rgba(0,0,0,.2);box-shadow:0px 10px 12px 5px rgba(0,0,0,.2)}.ndfHFb-c4YZDc-EglORb-haAclf .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c{margin:0 auto;transform:scale(1.7)}.ndfHFb-c4YZDc-EglORb-u0pjoe,.ndfHFb-c4YZDc-EglORb-ge6pde,.ndfHFb-c4YZDc-EglORb-Ujd07d{min-width:300px;position:absolute;text-align:center}.ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c{background-repeat:no-repeat;display:inline-block;height:19px;position:relative;top:3px;width:19px}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/v-spinner_dark.gif')!important}.ndfHFb-c4YZDc-e1YmVc.ndfHFb-c4YZDc .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/v-spinner_gray.gif')!important}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited){background-image:none!important;height:21px;width:21px;top:2px}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c .ndfHFb-aZ2wEe{display:block}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c .ndfHFb-vyDMJf-aZ2wEe{height:32px;width:32px;margin-left:-16px}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited){height:32px;width:32px}.ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS{font-size:19px;line-height:19px;margin-left:12px}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS{color:#1e1e1e}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS,.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS{display:none}.ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c{background-repeat:no-repeat;background-position:0 -800px;display:inline-block;height:37px;margin:0 auto;padding:0;width:31px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c{background-position:0 -2424px}.ndfHFb-c4YZDc-EglORb-u0pjoe-fmcmS,.ndfHFb-c4YZDc-EglORb-Ujd07d-fmcmS,.ndfHFb-c4YZDc-EglORb-u0pjoe-hSRGPd-haAclf{display:inline-block;font-size:19px;line-height:27px;-moz-user-select:text}.ndfHFb-c4YZDc-EglORb-Ujd07d-fmcmS{margin-top:15px}.ndfHFb-c4YZDc-EglORb-u0pjoe-hSRGPd-haAclf .ndfHFb-c4YZDc-EglORb-u0pjoe-KY1xSc-z5C9Gb-hSRGPd:link,.ndfHFb-c4YZDc-EglORb-u0pjoe-hSRGPd-haAclf .ndfHFb-c4YZDc-EglORb-u0pjoe-KY1xSc-z5C9Gb-hSRGPd:visited{padding-left:5px;color:#fff;cursor:pointer;display:inline-block;text-decoration:underline}.ndfHFb-c4YZDc-EglORb-u0pjoe-EbqdBd-ebJZBb-fmcmS{display:block;font-size:17px}.ndfHFb-c4YZDc-EglORb-u0pjoe-EbqdBd-ebJZBb{display:block;font-size:12px;text-align:left;white-space:pre-wrap;-moz-user-select:text}.ndfHFb-c4YZDc-EglORb-joDrKf-u0pjoe-fmcmS{font-size:13px;margin-top:10px}.ndfHFb-c4YZDc-EglORb-u0pjoe-Hr33Cd{font-size:19px;line-height:27px}.ndfHFb-c4YZDc-EglORb-nupQLb-LgbsSe,.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe{display:inline-block}.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe{margin-left:20px;margin-top:20px;-moz-border-radius:2px;border-radius:2px;background-color:#f5f5f5;background-image:-moz-linear-gradient(top,#f5f5f5,#f1f1f1);background-image:linear-gradient(top,#f5f5f5,#f1f1f1);border:1px solid #dcdcdc;border:1px solid rgba(0,0,0,.1);color:#444;font-size:11px;font-weight:bold;height:28px;line-height:28px;min-width:72px;outline:0;padding:0 8px;vertical-align:middle}.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe{-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1);background-color:#f8f8f8;background-image:-moz-linear-gradient(top,#f8f8f8,#f1f1f1);background-image:linear-gradient(top,#f8f8f8,#f1f1f1);border:1px solid #c6c6c6;color:#333}.ndfHFb-c4YZDc-LgbsSe-auswjd.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe{-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1);background-color:#f8f8f8;background-image:-moz-linear-gradient(top,#f8f8f8,#f1f1f1);background-image:linear-gradient(top,#f8f8f8,#f1f1f1);border:1px solid #c6c6c6;color:#333;-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.1);box-shadow:inset 0 1px 2px rgba(0,0,0,.1)}.ndfHFb-c4YZDc-LgbsSe-XpnDCe.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe{border:1px solid #4d90fe}.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe-Bz112c{background-size:contain;height:16px;left:10px;position:absolute;top:6px;width:16px}.ndfHFb-c4YZDc-EDpFhf-z5C9Gb-IyROMc-LgbsSe-fmcmS{margin-left:35px}.ndfHFb-c4YZDc-bN97Pc-u0pjoe-haAclf{color:#fff;padding-bottom:20px;text-align:center}.ndfHFb-c4YZDc-bN97Pc-u0pjoe-fmcmS{display:inline-block;font-size:15px;padding-left:20px;text-align:left;vertical-align:top}.XkWAb-LmsqOc{image-rendering:optimizeSpeed;image-rendering:-webkit-optimize-contrast;-moz-transition:opacity .5s linear;transition:opacity .5s linear}.XkWAb-xzdHvd{-moz-transform:translate(-50%,-50%) rotate(90deg) translate(50%,-50%);transform:translate(-50%,-50%) rotate(90deg) translate(50%,-50%)}.XkWAb-hTN0Jd{-moz-transform:translate(-50%,-50%) rotate(180deg) translate(-50%,-50%);transform:translate(-50%,-50%) rotate(180deg) translate(-50%,-50%)}.XkWAb-IZxJAe{-moz-transform:translate(-50%,-50%) rotate(270deg) translate(-50%,50%);transform:translate(-50%,-50%) rotate(270deg) translate(-50%,50%)}.XkWAb-cYRDff img.XkWAb-Iak2Lc{-moz-transition:none;transition:none}.XkWAb-cYRDff img.L6cTce{filter:alpha(opacity=0);opacity:0}.XkWAb-CHX6zb{filter:alpha(opacity=0);opacity:0;position:absolute;z-index:1002;height:100%;width:100%;background-color:#008000}.XkWAb-pfZwlb{overflow:hidden}.XkWAb-cYRDff{background:transparent!important;position:absolute;overflow:hidden}.XkWAb-LmsqOc{position:absolute}.XkWAb-pVNTue{position:absolute;z-index:1003;width:1px;height:1px;-moz-user-select:none}.XkWAb-RCfa3e{-moz-transition:all .5s;transition:all .5s}.XkWAb-pVNTue.XkWAb-RCfa3e{-moz-transition:opacity .5s;transition:opacity .5s}.XkWAb-pVNTue .XkWAb-sM5MNb{width:100%;height:100%;border:1px solid #808080;background:#000}.XkWAb-pVNTue .XkWAb-SMWX4b{direction:ltr;width:100%;height:100%;background-repeat:no-repeat;overflow:hidden;position:relative}.XkWAb-pVNTue .XkWAb-SMWX4b .XkWAb-pfZwlb .XkWAb-cYRDff{position:absolute}.XkWAb-pVNTue .XkWAb-xJ5Hz{background:transparent!important;border:1px solid #fff;position:absolute;z-index:1001}.XkWAb-pVNTue .XkWAb-ZdFRdf{position:absolute;background:#000;filter:alpha(opacity=60);opacity:.6;z-index:1001}.XkWAb-pVNTue .XkWAb-UH1Jve{width:100%;height:30px;background:#000;border-style:solid;border-color:#808080;border-width:0 1px 1px 1px;position:absolute;-moz-transition:height .5s;transition:height .5s}.XkWAb-eJuzjc,.XkWAb-a4WLyb{color:#fff;cursor:pointer;font-size:13px;height:30px;position:absolute;top:0;text-align:center;-moz-transition:height .5s;transition:height .5s;vertical-align:middle;width:22px}.XkWAb-BtWyge{display:table-cell;width:22px;height:30px;text-align:center;vertical-align:middle}.XkWAb-pVNTue .XkWAb-eJuzjc{right:0}.XkWAb-pVNTue .XkWAb-a4WLyb{left:0}.XkWAb-pVNTue .XkWAb-IlRY5e{height:30px;width:16px;background:#fff!important;cursor:pointer;-moz-transition:height .5s;transition:height .5s}.XkWAb-pVNTue .XkWAb-IE9qgd{left:22px;position:absolute;right:22px;top:0;-moz-transition:height .5s;transition:height .5s}.XkWAb-AHe6Kc{background-image:url("data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAACAAAAAgAQMAAABJtOi3AAAAAXNSR0IArs4c6QAAAAZQTFRF9/f3////TOsULwAAABRJREFUCNdjYGD4/5+BigR1TWMAAO29P8H0ss2LAAAAAElFTkSuQmCC");position:absolute;z-index:1}.ndfHFb-c4YZDc-ls4dqb{position:absolute;left:0;right:0;top:0;bottom:0;z-index:1}.XkWAb-cYRDff,.XkWAb-xJ5Hz{background-color:transparent!important}.XkWAb-pVNTue .XkWAb-IlRY5e{background-color:#fff!important}.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=87);opacity:0.87;background-position:0 -160px;margin-left:auto;margin-right:auto;margin-top:3px;height:21px;width:21px}.ndfHFb-c4YZDc-z5C9Gb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-z5C9Gb-LgbsSe-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -400px;margin-top:2px;height:24px;width:24px}.ndfHFb-c4YZDc-z5C9Gb-LgbsSe-ndfHFb-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -1920px;margin-top:2px;height:24px;width:24px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -2746px;margin-top:0;height:24px;width:24px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-z5C9Gb-LgbsSe-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -1568px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-z5C9Gb-LgbsSe-ndfHFb-yEEHq.ndfHFb-c4YZDc-z5C9Gb-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -328px}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-z5C9Gb-xl07Ob{font-size:13px;min-width:240px;padding:8px 0}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-Bz112c{filter:alpha(opacity=60);opacity:.6;left:12px;top:6px;margin-left:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-Bz112c{opacity:1}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c{top:5px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-j7LFlb-sn54Q .ndfHFb-c4YZDc-j7LFlb-Bz112c{top:6px}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-z5C9Gb-xl07Ob .ndfHFb-c4YZDc-z5C9Gb-xl07Ob-xl07Ob-ibnC6b-OWB6Me{filter:alpha(opacity=60);opacity:.6}.ndfHFb-c4YZDc-tJiF1e-LgbsSe,.ndfHFb-c4YZDc-E7ORLb-LgbsSe{position:absolute;top:80px;bottom:80px;margin-top:auto;margin-bottom:auto;outline:0;width:40px;height:90px;z-index:5}.ndfHFb-c4YZDc-tJiF1e-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-E7ORLb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-tJiF1e-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -1960px}.ndfHFb-c4YZDc-E7ORLb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -840px}.ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -1640px}.ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -680px}.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c:not([onclick]):not(:link):not(:visited),.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url(//ssl.gstatic.com/docs/common/v-icons4.png)!important}.ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:-26px -26px}.ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -248px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -2096px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -248px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe.ndfHFb-c4YZDc-PRu6Hd-QebRhd.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -2096px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tJiF1e-LgbsSe,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-E7ORLb-LgbsSe{width:48px}.ndfHFb-c4YZDc-DH6Rkf-Bz112c{height:24px;position:absolute;width:24px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-Bz112c{height:24px;width:24px}.ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{height:30px;width:40px;background:#000;-moz-border-radius:3px;border-radius:3px;filter:alpha(opacity=80);opacity:.8;position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{height:40px;width:40px;-moz-border-radius:20px;border-radius:20px;background:rgba(0,0,0,.75);-moz-transition:background 0.2s,opacity 0.34s,transform 0.34s cubic-bezier(0.4,0.0,0.2,1);transition:background 0.2s,opacity 0.34s,transform 0.34s cubic-bezier(0.4,0.0,0.2,1);opacity:1}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{background:var(--dt-surface,#fff)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc .ndfHFb-c4YZDc-DH6Rkf-Bz112c{position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{background:#4285f4}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{background:#696b6a}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-auswjd .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{background:#6d6f6f}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-LgbsSe-XpnDCe .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{outline:#4d90fe solid 1px}.ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-DH6Rkf-AHe6Kc{display:none}.ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d{display:inline-block;margin-right:10px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d{border:1px solid transparent;-moz-border-radius:2px;border-radius:2px;background:rgba(0,0,0,.75);margin:0;white-space:nowrap}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d{-moz-border-radius:100px;border-radius:100px;border-color:var(--dt-outline,#80868b);background-color:var(--dt-surface,#fff)}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe.ndfHFb-c4YZDc-Wrql6b-FNFY6c-BP2Omd-qMHh7d,.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c.ndfHFb-c4YZDc-Wrql6b-FNFY6c-BP2Omd-qMHh7d{border-bottom-right-radius:0;border-right:0;border-top-right-radius:0;display:inline-block;margin-right:0;min-width:64px}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c,.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d{font-size:13px;font-weight:normal;margin:0}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d{font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d{min-width:0;padding:0;color:white;height:30px;margin-left:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d{color:var(--dt-on-surface-variant,#5f6368);height:36px}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c{padding-right:4px;min-width:79px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c{padding-left:8px;padding-right:8px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-FNFY6c{padding-left:16px;padding-right:16px}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d{display:inline-block;min-width:89px;padding:10px 0}.ndfHFb-c4YZDc-FNFY6c-V67aGc{display:inline-block}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-V67aGc{line-height:24px;margin-top:4px;max-width:200px;overflow:hidden;text-overflow:ellipsis}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-V67aGc{margin-top:6px;margin-left:4px}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-Wrql6b-qMHh7d.ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp{border-bottom-left-radius:0;border-left:0;border-top-left-radius:0;min-width:15px}.ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS{display:inline-block;min-width:59px;padding-left:4px;padding-right:6px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS{line-height:30px;padding-left:8px;padding-right:0;float:left}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS{line-height:24px;padding-left:16px;padding-right:0;float:left;margin-top:4px}.ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS{display:none}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-Wrql6b-PlOyMe,.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-Wrql6b-FNFY6c,.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-Wrql6b-qMHh7d{background-color:#232323;background-image:-moz-linear-gradient(top,#333,#222);background-image:linear-gradient(top,#333,#222)}.ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb,.ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb{display:inline-block;margin:0 4px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb{margin:0;overflow:hidden}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb{margin-top:2px}.ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo{filter:alpha(opacity=80);opacity:.8;display:inline-block;margin-bottom:1px;vertical-align:middle}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo{filter:alpha(opacity=100);opacity:1;border-bottom-right-radius:2px;border-right:2px;border-top-right-radius:2px;margin-bottom:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo{width:20px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:center;padding-right:12px;padding-left:4px}.ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo .ndfHFb-c4YZDc-Bz112c{background-position:0 -960px;height:16px;width:16px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo .ndfHFb-c4YZDc-Bz112c{background-position:0 -1936px;height:24px;width:24px;margin-top:4px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo .ndfHFb-c4YZDc-Bz112c{height:20px;width:20px}.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c{background-size:contain;display:inline-block;height:16px;margin-right:6px;width:16px;vertical-align:text-bottom}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c{float:left;height:24px;width:24px;margin-top:4px;margin-left:-4px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c{height:14px;width:14px;margin-top:11px;margin-bottom:11px;margin-left:2px}.ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe{border-left:1px solid rgba(255,255,255,.3);display:inline-block;height:11px;vertical-align:middle}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe{border-color:rgba(255,255,255,.35);height:24px;margin-top:3px;vertical-align:top}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-qMHh7d-yolsp .ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe{border-color:var(--dt-outline,#80868b);height:36px;width:1px;margin-top:0}.ndfHFb-c4YZDc-LgbsSe-ZmdkE~.ndfHFb-c4YZDc-Wrql6b-qMHh7d>.ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe,.ndfHFb-c4YZDc-LgbsSe-ZmdkE>.ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe{opacity:0}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe-ZmdkE~.ndfHFb-c4YZDc-Wrql6b-qMHh7d>.ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe-ZmdkE>.ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe{opacity:100%}.ndfHFb-c4YZDc-DARUcf-NnAfwf{-moz-transition:opacity .218s;transition:opacity .218s;background-color:#000;-moz-border-radius:3px;border-radius:3px;bottom:10px;position:absolute;line-height:25px;padding:0 18px;text-align:center;height:25px;min-width:56px;z-index:3}.ndfHFb-c4YZDc-DARUcf-NnAfwf-auswjd{filter:alpha(opacity=70);opacity:.7}.ndfHFb-c4YZDc-DARUcf-NnAfwf-L6cTce{filter:alpha(opacity=0);opacity:0}.ndfHFb-c4YZDc-DARUcf-NnAfwf-fmcmS{color:#fff;font-size:11px;font-weight:bold}.ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb{border-right:1px solid rgba(255,255,255,.2);display:inline-block;font-size:13px;line-height:44px;height:44px;vertical-align:middle}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em);display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center}.ndfHFb-c4YZDc-DARUcf-NnAfwf-tJHJj{display:inline-block;margin-left:12px;vertical-align:middle}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-DARUcf-NnAfwf-tJHJj{margin-left:16px}.ndfHFb-c4YZDc-DARUcf-NnAfwf-cQYSPc,.ndfHFb-c4YZDc-DARUcf-NnAfwf-j4LONd{display:inline-block;text-align:center;vertical-align:middle;width:48px}.ndfHFb-c4YZDc-cYSp0e,.ndfHFb-c4YZDc-cYSp0e-s2gQvd{bottom:0;left:0;position:absolute;right:0;top:0}.ndfHFb-c4YZDc-cYSp0e-Oz6c3e{position:relative}.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e{max-width:800px;margin-left:auto;margin-right:auto;margin-top:60px;margin-bottom:60px}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e{margin-top:56px;margin-bottom:56px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e{margin-top:64px;margin-bottom:64px}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-TJEFFc.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-cYSp0e-Oz6c3e{margin-top:12px;margin-bottom:12px}.ndfHFb-c4YZDc-cYSp0e-hpYHOb{bottom:0;position:absolute;top:0}.ndfHFb-c4YZDc-cYSp0e{outline:none}.ndfHFb-c4YZDc-cYSp0e-BIzmGd{border:1px solid #eee;-moz-box-shadow:0 3px 3px rgba(0,0,0,.05);box-shadow:0 3px 3px rgba(0,0,0,.05);background:rgba(255,255,255,.95);-moz-border-radius:100%;border-radius:100%;display:block;opacity:0;position:absolute;width:40px;height:40px;left:100%;margin-left:-22px;cursor:pointer;transition:opacity .25s ease-in-out;z-index:3}.ndfHFb-c4YZDc-cYSp0e-BIzmGd.ndfHFb-c4YZDc-LgbsSe{opacity:1}.ndfHFb-c4YZDc-cYSp0e-BIzmGd.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me{opacity:0}.ndfHFb-c4YZDc-BIzmGd-Bz112c{background-position:0 -2642px;display:inline-block;height:24px;margin:10px 10px;opacity:.5;pointer-events:none;width:24px}.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-cYSp0e-BIzmGd .ndfHFb-c4YZDc-BIzmGd-Bz112c{opacity:1}.ndfHFb-c4YZDc-cYSp0e-s2gQvd{overflow:auto}.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-s2gQvd{margin-left:12px;margin-right:12px;overflow:hidden}.ndfHFb-c4YZDc-cYSp0e-B7I4Od{left:-5000px;position:absolute;top:-5000px}.ndfHFb-c4YZDc-cYSp0e-DARUcf{position:relative;pointer-events:none;background-color:rgba(79,79,79,.2)}.ndfHFb-c4YZDc-cYSp0e-DARUcf+.ndfHFb-c4YZDc-cYSp0e-DARUcf{margin-top:40px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-cYSp0e-DARUcf+.ndfHFb-c4YZDc-cYSp0e-DARUcf{margin-top:16px}.ndfHFb-c4YZDc.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-cYSp0e-DARUcf+.ndfHFb-c4YZDc-cYSp0e-DARUcf{margin-top:12px}.ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf{font-size:11px;opacity:.01;overflow:hidden;height:100%;position:absolute;width:100%;z-index:-1}.ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj,.ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe{position:absolute;margin:0;padding:0;border-width:0}.ndfHFb-c4YZDc-cYSp0e-DARUcf-gSKZZ .ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf{cursor:text}.ndfHFb-c4YZDc-cYSp0e-DARUcf-xUXeUb .ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf{cursor:crosshair}.ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c{position:absolute;width:100%;height:100%;-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35)}.ndfHFb-c4YZDc-cYSp0e-DARUcf-M1R4Ee-UzWXSb{position:absolute;width:100%;height:100%;-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);background-color:#fff}.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c{-moz-box-shadow:none;box-shadow:none}.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-DARUcf{background-color:transparent}.ndfHFb-c4YZDc-TJEFFc .ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c{position:relative;height:auto}.ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf{height:100%;overflow:hidden;position:absolute;width:100%;pointer-events:auto;z-index:2}.ndfHFb-c4YZDc-cYSp0e-DARUcf-hSRGPd{cursor:pointer;position:absolute;background-image:url(data:image/gif;base64,R0lGODlhAQABAIAAAP///wAAACH5BAEAAAAALAAAAAABAAEAAAICRAEAOw==)}.ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q{position:absolute;filter:alpha(opacity=35);opacity:.35;background-color:#ffe168;z-index:1}.ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-bN97Pc-u0pjoe-haAclf,.ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-EglORb-ge6pde{position:relative}.ndfHFb-c4YZDc-cYSp0e-DARUcf-u0pjoe-DARUcf{position:absolute;height:100%;width:100%;pointer-events:auto;z-index:2}.ndfHFb-c4YZDc-cYSp0e-DARUcf-u0pjoe-EglORb{text-align:center;width:100%;position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-bN97Pc-u0pjoe-fmcmS{font-size:15px;line-height:25px}.ndfHFb-c4YZDc-cYSp0e .ndfHFb-c4YZDc-EglORb-u0pjoe-RJLb9c{margin:5px 0}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf:not([onclick]):not(:link):not(:visited){background-color:transparent!important}.ndfHFb-c4YZDc-UmsTj-Sx9Kwc{position:absolute;min-width:400px;height:105px;background:#232323;border:1px solid #000;-moz-border-radius:3px;border-radius:3px;color:white;cursor:default;font-size:15px;font-weight:bold;font-family:arial,sans-serif;-moz-user-select:text}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Sx9Kwc{background:var(--dt-surface,#fff);padding:24px 24px;-moz-border-radius:8px;border-radius:8px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center;flex-direction:column;justify-content:space-between;height:auto}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Sx9Kwc-ma6Yeb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;margin:0 0 24px 0}.ndfHFb-c4YZDc-UmsTj-Ne3sFf{position:relative;top:11px;margin-left:40px;margin-right:10px;white-space:nowrap}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Ne3sFf{position:static;font:var(--dt-title-large-font,400 1.375rem/1.75rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-title-large-spacing,0);margin:0 16px}.ndfHFb-c4YZDc-UmsTj-Bz112c{position:absolute;top:4px;left:7px;width:28px;height:28px;background-position:0 -920px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UmsTj-Bz112c{background-position:0 -1328px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UmsTj-Bz112c{background-position:0 -472px;position:static}.ndfHFb-c4YZDc-UmsTj-YPqjbf-sM5MNb{position:absolute;left:10px;right:10px;top:40px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-YPqjbf-sM5MNb{position:static;width:100%}.ndfHFb-c4YZDc-UmsTj-YPqjbf{position:absolute;top:0;height:19px;width:100%;margin:0;background-color:#5c5c5c;border:1px solid #000;color:white;font:normal 16px arial,sans-serif;box-sizing:content-box;-moz-box-sizing:content-box}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-YPqjbf{position:static;height:26px;box-sizing:border-box}.ndfHFb-c4YZDc-UmsTj-Sx9Kwc-cGMI2b{position:relative;top:53px;width:100%;white-space:nowrap}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-Sx9Kwc-cGMI2b{position:static;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;justify-content:space-between;margin:24px 0 0 0}.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf{top:0;right:9px;background-color:#4d90fe;color:rgba(255,255,255,.87);margin:0;padding:0 8px;font-size:13px;height:25px;line-height:25px;min-width:50px;text-align:center}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf{-moz-border-radius:100px;border-radius:100px;background:var(--dt-surface,#fff);color:var(--dt-primary,#1a73e8);font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em);border:none;margin:0;padding:0;position:static;height:30px;min-width:72px;line-height:30px}.ndfHFb-c4YZDc-UmsTj-u0pjoe{top:2px;min-width:295px;white-space:nowrap;display:inline-block;position:static;margin:0}.ndfHFb-c4YZDc-UmsTj-u0pjoe-fmcmS{color:#f00}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-UmsTj-u0pjoe-fmcmS{color:var(--dt-error,#d93025);font:var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-large-spacing,0.00625em);height:30px;line-height:30px}.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me.ndfHFb-c4YZDc-UmsTj-sFeBqf{background-color:#808080;color:#c2c2c2}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me.ndfHFb-c4YZDc-UmsTj-sFeBqf{background:var(--dt-surface,#fff);color:var(--dt-on-surface,#3c4043);opacity:.38}.ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-UmsTj-sFeBqf{background-color:#4d90fe;background-image:-moz-linear-gradient(top,#4d90fe,#357ae8);background-image:linear-gradient(top,#4d90fe,#357ae8);color:rgba(255,255,255,1)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-UmsTj-sFeBqf{background:rgba(168,199,250,.08);color:var(--dt-primary,#1a73e8);border:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf:focus,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-UmsTj-sFeBqf:active{background:rgba(168,199,250,.12);color:var(--dt-primary,#1a73e8);border:none;outline:none;-moz-box-shadow:none;box-shadow:none}.ndfHFb-c4YZDc-n1UuX-Bz112c,.ndfHFb-c4YZDc-mKZypf-bEDTcc,.ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-yHKmmc,.ndfHFb-c4YZDc-no16zc-UcSZ6e{display:inline-block;padding:9px 0}.ndfHFb-c4YZDc-Woal0c-jcJzye-ZMv3u{vertical-align:middle}.ndfHFb-c4YZDc-n1UuX-RJLb9c{background-color:#464445;-moz-border-radius:50%;border-radius:50%;height:29px;width:29px;margin-left:13px;vertical-align:middle}.ndfHFb-c4YZDc-no16zc-UcSZ6e{vertical-align:middle}.ndfHFb-c4YZDc-no16zc-UcSZ6e-LgbsSe{margin-left:13px;margin-right:0;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.ndfHFb-c4YZDc-mKZypf-bEDTcc-LgbsSe{margin-left:13px;margin-right:0}.ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-LgbsSe,.ndfHFb-c4YZDc-UcSZ6e-mKZypf-yHKmmc-LgbsSe{display:inline-block;margin-left:13px;margin-right:0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-n1UuX-Bz112c{padding:5.5px 8px 5.5px 8px;margin-left:3px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-mKZypf-bEDTcc,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-yHKmmc,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-no16zc-UcSZ6e{padding:5.5px 8px 5.5px 8px;margin-left:8px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-n1UuX-RJLb9c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-mKZypf-bEDTcc-LgbsSe,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-no16zc-UcSZ6e-LgbsSe,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-LgbsSe,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-yHKmmc-LgbsSe{margin-left:0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-UcSZ6e-mKZypf-bEDTcc-LgbsSe+.ndfHFb-c4YZDc-UcSZ6e-mKZypf-yHKmmc-LgbsSe{margin-left:13px}.ndfHFb-c4YZDc-kODWGd-umzg3c{height:100%;position:absolute;left:46px;right:auto}.ndfHFb-c4YZDc-kODWGd-umzg3c-SxecR{width:130px}.ndfHFb-c4YZDc-kODWGd-umzg3c-SxecR-PFprWc{height:12px;width:20px}.ndfHFb-c4YZDc-kODWGd-umzg3c-ihIZgd{font-family:"Open Sans",arial,sans-serif;font-size:13px;font-weight:bold;min-width:30px;top:8px;left:144px;right:auto;position:absolute}.ndfHFb-c4YZDc-sbW6Cb{-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);background-color:#f8f8f8;color:#2a2a2a;display:block;font:13px "Google Sans",arial,sans-serif;line-height:19px;margin-left:20px;opacity:1;position:absolute;visibility:visible;z-index:1294}.ndfHFb-c4YZDc-sbW6Cb-bN97Pc{padding:10px}.ndfHFb-c4YZDc-sbW6Cb-bN97Pc-hSRGPd{color:#2a2a2a;text-decoration:underline}.ndfHFb-c4YZDc-sbW6Cb-hFsbo{position:absolute}.ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe,.ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{content:"";display:block;height:0;position:absolute;width:0}.ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe{border:16px solid}.ndfHFb-c4YZDc-sbW6Cb-hFsbo .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{border:14px solid}.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb{bottom:0}.ndfHFb-c4YZDc-sbW6Cb-d6mlqf{top:-14px}.ndfHFb-c4YZDc-sbW6Cb-y6n2Me{left:-14px}.ndfHFb-c4YZDc-sbW6Cb-cX0Lwc{right:0}.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe,.ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe{border-color:#f8f8f8 transparent;left:-16px}.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc,.ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{border-color:#f8f8f8 transparent;left:-14px}.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe,.ndfHFb-c4YZDc-sbW6Cb-Ya1KTb .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{border-bottom-width:0}.ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe{border-top-width:0}.ndfHFb-c4YZDc-sbW6Cb-d6mlqf .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{border-top-width:0;top:2px}.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe,.ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe{border-color:transparent #f8f8f8;top:-16px}.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc,.ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{border-color:transparent #f8f8f8;top:-14px}.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe{border-left-width:0}.ndfHFb-c4YZDc-sbW6Cb-y6n2Me .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{border-left-width:0;left:2px}.ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-WgXLxe,.ndfHFb-c4YZDc-sbW6Cb-cX0Lwc .ndfHFb-c4YZDc-sbW6Cb-Zj4Smb-BuvAkc{border-right-width:0}.ndfHFb-c4YZDc-Lo93Wb-fmcmS{display:inline-block;vertical-align:middle;max-width:150px;margin-right:5px}.ndfHFb-c4YZDc-Lo93Wb-Bz112c{display:inline-block;vertical-align:middle;background-repeat:no-repeat;filter:alpha(opacity=87);opacity:0.87;height:21px;width:21px}.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc{color:#000;font:normal 13px arial,sans-serif;width:340px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc{color:var(--dt-on-surface,#3c4043);font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-r4nke{font-weight:normal;margin:0 0 16px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-r4nke{margin:0 0 24px}.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc{-moz-border-radius:1px;border-radius:1px;border:1px solid #d9d9d9;border-top:1px solid #c0c0c0;font-size:13px;height:25px;padding:1px 8px;width:300px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc{border:2px solid var(--dt-primary,#1a73e8);font:var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-large-spacing,0.00625em);padding:8px 16px;-moz-border-radius:4px;border-radius:4px;background:var(--dt-surface,#fff);color:var(--dt-on-surface,#3c4043)}.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc:focus{-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.3);box-shadow:inset 0 1px 2px rgba(0,0,0,.3);border:1px solid #4d90fe;outline:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc:focus{border:2px solid var(--dt-primary,#1a73e8)}.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-dI4VCc::-ms-clear{display:none}.ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-c6xFrd{margin-top:16px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-c6xFrd{margin-top:24px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:flex-end}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Iqlsrf-Sx9Kwc-c6xFrd button{cursor:pointer}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Iqlsrf-Bz112c{background-position:0 -976px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Iqlsrf-Bz112c{background-position:0 -856px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Sx9Kwc-bN97Pc br{display:none}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe{position:absolute;left:-300px;top:-42px;z-index:4;height:40px;width:295px;background-color:#2d2d2d;border:1px solid #000;-moz-border-radius:3px;border-radius:3px;border-top-width:1px;-moz-transition:top .218s ease-out;transition:top .218s ease-out}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe{left:-600px;background:var(--dt-surface3,#fff);-moz-box-shadow:0 4px 8px 3px rgba(0,0,0,.15),0 1px 3px rgba(0,0,0,.3);box-shadow:0 4px 8px 3px rgba(0,0,0,.15),0 1px 3px rgba(0,0,0,.3);-moz-border-radius:8px;border-radius:8px;padding:12px 16px;border:none;height:36px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center;width:336px}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-ti6hGc,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-ti6hGc{left:unset;right:56px;top:50px}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf{position:relative;margin:0 0 0 4px;vertical-align:middle;height:25px;padding:0 9px;width:198px;background-color:#0a0a0a;border:solid #444;border-width:0 0 1px 1px;display:inline-block}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center;width:200px;height:auto;margin:0;padding:4px 8px;background:var(--dt-surface3,#fff);border:1px solid var(--dt-outline,#80868b);-moz-border-radius:4px;border-radius:4px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf:hover{border:1px solid var(--dt-on-surface,#3c4043)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf-XpnDCe{border:2px solid var(--dt-primary,#1a73e8)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf-x5ghY{border:2px solid var(--dt-error,#d93025)}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf-haAclf{display:table-cell;width:100%}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf,.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf{color:#fff;font-size:13px;font-weight:normal}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf{width:100%;background-color:#0a0a0a;border:0;height:25px;outline:none!important;padding:0}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf{height:24px;font:var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-large-spacing,0.00625em);background:var(--dt-surface3,#fff)}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf::-webkit-input-placeholder{color:#fff;opacity:.75}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf::-moz-placeholder{color:#fff;opacity:.75}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf:-ms-input-placeholder{color:#fff;opacity:.75}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf-haAclf{display:table-cell;max-width:100px;opacity:.5;padding-left:7px;white-space:nowrap}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf{padding:0 2px}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf-x5ghY{background-color:#ff4500}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne{position:relative;top:8px;height:21px;width:21px;opacity:.7}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne{position:static;top:0;opacity:1;-moz-border-radius:100px;border-radius:100px;margin-left:8px;padding:8px;height:21px;width:21px}.ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne{opacity:.9}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-LgbsSe-ZmdkE.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne{opacity:1}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:rgba(196,199,197,.08)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-LgbsSe-XpnDCe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-LgbsSe-auswjd{background-color:rgba(196,199,197,.12)}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc{background-position:0 0;margin-left:-2px;top:5px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc{top:0;margin-left:8px;height:21px;width:21px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc .ndfHFb-c4YZDc-Bz112c{transform:scale(0.86);position:relative;top:-1px;right:1px}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc.ndfHFb-c4YZDc-w5vlXd{top:8px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc.ndfHFb-c4YZDc-w5vlXd{top:-1px}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e,.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb{border:1px solid #444}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb{border:none}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e{background-position:0 -80px;left:-1px;border-top-right-radius:3px;border-bottom-right-radius:3px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e .ndfHFb-c4YZDc-Bz112c{position:relative;top:1px}.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb{background-position:0 -1240px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc{background-position:0 -3178px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e{background-position:0 -1752px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb{background-position:0 -3754px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne .ndfHFb-c4YZDc-Bz112c{height:21px;width:21px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne.ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc .ndfHFb-c4YZDc-Bz112c{background-position:0 -3178px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e .ndfHFb-c4YZDc-Bz112c{background-position:0 -1752px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb .ndfHFb-c4YZDc-Bz112c{background-position:0 -3754px}.ndfHFb-c4YZDc-O1htCb-LgbsSe,.ndfHFb-c4YZDc-O1htCb-K2kob{background-color:rgba(90,90,90,.7);border:2px solid #d7d7d7;height:32px;left:70px;position:absolute;top:80px;width:32px;z-index:5;-moz-border-radius:50%;border-radius:50%}@media screen and (max-width:800px){.ndfHFb-c4YZDc-O1htCb-LgbsSe{left:5%}}.ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE,.VIpgJd-j7LFlb-sn54Q .ndfHFb-c4YZDc-O1htCb-K2kob{background-color:rgba(138,138,138,.7);border:2px solid #fff;-moz-box-shadow:0px 2px 5px rgba(83,83,83,.7);box-shadow:0px 2px 5px rgba(83,83,83,.7)}.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-O1htCb-LgbsSe,.VIpgJd-wQNmvb-gk6SMd .ndfHFb-c4YZDc-O1htCb-K2kob{background-color:#4d90fe;border:2px solid #fff;-moz-box-shadow:0px 2px 5px rgba(83,83,83,.7);box-shadow:0px 2px 5px rgba(83,83,83,.7)}.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE,.VIpgJd-wQNmvb-gk6SMd.VIpgJd-j7LFlb-sn54Q .ndfHFb-c4YZDc-O1htCb-K2kob{background-color:#5e9bfe}.ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-O1htCb-LgbsSe-gk6SMd-YLEHIf,.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b-YLEHIf .ndfHFb-c4YZDc-O1htCb-K2kob{-moz-animation:driveViewerSelectButtonSelectedAnimation .3s linear 0s 1;animation:driveViewerSelectButtonSelectedAnimation .3s linear 0s 1}.ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c,.ndfHFb-c4YZDc-O1htCb-K2kob-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v-sprite19.svg');background-position:0 -1320px;width:30px;height:30px;margin-top:-4px;filter:alpha(opacity=70);opacity:.7}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c,.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-O1htCb-K2kob-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -2682px}.ndfHFb-c4YZDc-O1htCb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c{filter:alpha(opacity=90);opacity:.9}.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-O1htCb-LgbsSe-Bz112c{filter:alpha(opacity=100);opacity:1}@-moz-keyframes driveViewerSelectButtonSelectedAnimation{0%{opacity:.3}50%{opacity:1}}@keyframes driveViewerSelectButtonSelectedAnimation{0%{opacity:.3}50%{opacity:1}}.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob{background:#ededed;-moz-border-radius:3px;border-radius:3px;border:none;-moz-box-shadow:0 1px 2px 1px rgba(0,0,0,.4);box-shadow:0 1px 2px 1px rgba(0,0,0,.4);margin-top:4px;margin-left:-35px;max-height:70%;max-width:645px}.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-j7LFlb{display:inline-block;padding:0}.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-j7LFlb-sn54Q{padding:0;border:none}.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-JUCs7e{border:none;-moz-border-radius:0;border-radius:0;display:block;height:auto;margin:0;width:auto}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b{display:inline-block;height:110px;margin:3px 8px;overflow:hidden;position:relative;width:110px}.ndfHFb-c4YZDc-gvZm2b-xl07Ob .ndfHFb-c4YZDc-JUCs7e-SmKAyb{display:table-cell;height:90px;text-align:center;vertical-align:middle;width:110px}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-JUCs7e-SmKAyb img{-moz-box-shadow:0 1px 2px 0 rgba(0,0,0,.7);box-shadow:0 1px 2px 0 rgba(0,0,0,.7);max-width:100%;max-height:90%;display:inline-block}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b img.ndfHFb-c4YZDc-JUCs7e-Bz112c{background-color:#f5f5f5;height:60px;width:60px}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b-r4nke{font-size:15px;margin-top:3px;overflow:hidden;text-overflow:ellipsis;text-align:center;white-space:nowrap}@media screen and (max-width:1350px){.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob{max-width:520px}}@media screen and (max-width:1000px){.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob{max-width:390px}}@media screen and (max-width:700px){.ndfHFb-c4YZDc-xl07Ob.ndfHFb-c4YZDc-gvZm2b-xl07Ob{max-width:273px}}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob-Bz112c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob{position:absolute;right:0;top:55px}.VIpgJd-j7LFlb-sn54Q .ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob,.VIpgJd-wQNmvb-gk6SMd .ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b .ndfHFb-c4YZDc-O1htCb-K2kob{-moz-box-shadow:none;box-shadow:none}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.VIpgJd-wQNmvb-gk6SMd{background-image:none}.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.VIpgJd-j7LFlb-sn54Q,.ndfHFb-c4YZDc-gvZm2b-xl07Ob-ibnC6b.VIpgJd-j7LFlb-ZmdkE{background-color:transparent;border:none;padding:0}.ndfHFb-c4YZDc-uoC0bf .euCgFf-X3SwIb-haAclf{padding:0}.ndfHFb-c4YZDc-ZCZpd-h9d3hd{-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);outline:none;z-index:1293!important}.ndfHFb-c4YZDc-qbOKL-OEVmcd .IyROMc-w3KqTd-ztA2jd-SUR3Rd{z-index:1294!important}.ndfHFb-c4YZDc-SxecR{height:12px;margin-top:12px;padding-left:0;padding-right:2px}.ndfHFb-c4YZDc-SxecR-PFprWc{background-color:#e5e5e5;background-image:-moz-linear-gradient(top,#fff,#c0c0c0);background-image:linear-gradient(top,#fff,#c0c0c0);-moz-box-shadow:0 0 5px 0px #000;box-shadow:0 0 5px 0px #000;background-color:#e5e5e5!important;-moz-border-radius:6px;border-radius:6px;position:absolute;top:10px}.ndfHFb-c4YZDc-SxecR-skjTt{-moz-border-radius:8px;border-radius:8px;height:6px;position:absolute}.ndfHFb-c4YZDc-SxecR-cQwEuf{background-color:#4d4d4d;margin-top:1px;width:0}.ndfHFb-c4YZDc-SxecR-skjTt-j4LONd{background-color:transparent;border:1px solid #808080!important;width:inherit}.ndfHFb-c4YZDc-SxecR-skjTt-MFS4be{background-color:#d9d9d9;background-image:-moz-linear-gradient(top,#c3c3c3,#d9d9d9);background-image:linear-gradient(top,#c3c3c3,#d9d9d9);background-color:#d9d9d9!important;border-bottom-right-radius:0;border-top-right-radius:0;margin-top:1px;width:0}.ndfHFb-c4YZDc-Ng57nc.ndfHFb-c4YZDc-b3rLgd-haAclf{bottom:24px;left:24px;position:absolute;text-align:left;z-index:4}.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-Ng57nc.ndfHFb-c4YZDc-b3rLgd-haAclf{bottom:0;left:0;text-align:center;width:100%}.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd{-moz-border-radius:2px;border-radius:2px;-moz-box-shadow:0px 2px 4px rgba(0,0,0,.2);box-shadow:0px 2px 4px rgba(0,0,0,.2);align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-transform:translate3d(0,72px,0);transform:translate3d(0,72px,0);-moz-transition:transform .15s cubic-bezier(0.4,0.0,1,1),opacity .15s cubic-bezier(0.4,0.0,1,1),visibility 0ms linear .15s;transition:transform .15s cubic-bezier(0.4,0.0,1,1),opacity .15s cubic-bezier(0.4,0.0,1,1),visibility 0ms linear .15s;-moz-transition:all 0 linear 1s,opacity 1s;transition:all 0 linear 1s,opacity 1s;background-color:#eee;border:none;color:black;font-size:14px;margin:0;max-width:568px;min-height:20px;min-width:288px;opacity:0;padding:14px 0 14px 24px;text-align:left}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd{background:var(--dt-surface,#fff);color:var(--dt-on-surface,#3c4043);padding:14px 8px 14px 24px}.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd{background-color:#323232;color:white;max-width:none;width:100%}.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-TSZdd{-moz-transition-delay:0s;transition-delay:0s;-moz-transform:translate3d(0,0,0);transform:translate3d(0,0,0);bottom:24px;opacity:1}.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-Ne3sFf{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;-moz-flex:1 1 0;flex:1 1 0;line-height:19px;overflow:hidden}.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd{-moz-flex:0 0 auto;flex:0 0 auto;padding-left:24px;padding-right:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd{text-transform:none;-moz-border-radius:100px;border-radius:100px;height:30px;line-height:30px;margin:0 8px 0 16px;padding:0 16px}.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd,.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd,.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited,.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:visited{background:none;border:none;color:#1967d2;cursor:pointer;font-family:inherit;font-size:inherit;font-weight:bold;margin:0;outline:none;text-decoration:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:visited{color:var(--dt-primary,#1a73e8)}.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd,.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:visited{text-transform:uppercase;float:right}.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover,.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:focus,.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:hover,.ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:focus{text-decoration:underline}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:focus,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:hover,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-hSRGPd:focus{text-decoration:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:hover{background:rgba(168,199,250,.08)}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:focus,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd:active{background:rgba(168,199,250,.12)}.ndfHFb-c4YZDc-N4imRe .ndfHFb-c4YZDc-Ng57nc .ndfHFb-c4YZDc-b3rLgd-JIbuQc-hSRGPd{color:#a1c2fa;padding-right:48px}.ndfHFb-c4YZDc-L7w45e-ORHb{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;background-color:#f9ab00;-moz-border-radius:0;border-radius:0;color:#202124;height:3rem;position:relative;top:0;width:100%;z-index:3}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb{background:#ffdf99}.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;background-color:var(--dt-error,#d93025);-moz-border-radius:0;border-radius:0;color:#fff;height:3rem;position:relative;top:0;width:100%;z-index:3}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb{background:#ec928e;color:#202124}.ndfHFb-c4YZDc-L7w45e-ORHb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3098px;height:24px;margin:0 25px;width:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-Bz112c{margin:0 16px}.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3714px;height:24px;margin:0 25px;width:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Bz112c{background-position:0 -3098px;margin:0 16px}.ndfHFb-c4YZDc-L7w45e-ORHb-bN97Pc,.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-bN97Pc{align-items:center;display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;justify-content:space-between;width:100%}.ndfHFb-c4YZDc-L7w45e-ORHb-Ne3sFf,.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Ne3sFf{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-Ne3sFf,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-Ne3sFf{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-L7w45e-ORHb-LQLjdd,.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-LQLjdd{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;align-items:center;margin:8px 0;-moz-box-ordinal-group:0;order:0}.ndfHFb-c4YZDc-L7w45e-ORHb-IYtByb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3570px}.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -3178px}.ndfHFb-c4YZDc-L7w45e-ORHb-IYtByb-Bz112c,.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-Bz112c{margin:0 16px;height:20px;width:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-IYtByb-Bz112c{background-position:0 -3570px}.ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe{align-self:center;color:#202124;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px;padding:4px 18px;text-align:center;text-decoration:none;-moz-border-radius:20px;border-radius:20px;border:1px solid black;border-color:black}.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe{align-self:center;color:#fff;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px;padding:4px 18px;text-align:center;text-decoration:none;-moz-border-radius:20px;border-radius:20px;border:1px solid white;border-color:white}.ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe{align-self:center;color:#202124;font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;letter-spacing:.25px;line-height:20px;padding:0 16px;text-align:center;text-decoration:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe{border:none;color:#202124;font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em);padding:0 12px;min-width:70px}.ndfHFb-c4YZDc-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe:hover,.ndfHFb-c4YZDc-L7w45e-ORHb-Rsbfue-LPmGke-LgbsSe:hover,.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb-JLm1tf-L7w45e-LgbsSe:hover{cursor:pointer}.ndfHFb-c4YZDc-L7w45e-ORHb.ndfHFb-c4YZDc-ORHb-L6cTce,.ndfHFb-c4YZDc-oKM7Re-L7w45e-ORHb.ndfHFb-c4YZDc-ORHb-L6cTce{display:none}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc{align-items:flex-start;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;padding:0;outline:none;position:absolute;width:468px;background:#fff;-moz-box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);box-shadow:0px 1px 3px 0px rgba(60,64,67,.30),0px 4px 8px 3px rgba(60,64,67,.15);-moz-border-radius:8px;border-radius:8px;z-index:1194}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc{background:var(--dt-surface,#fff);padding:24px 24px;-moz-border-radius:8px;border-radius:8px}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-xJ5Hnf{background-color:#000;height:100%;left:0;position:fixed;top:0;width:100%;z-index:1194}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-bN97Pc{color:#f1f3f4;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:column;justify-content:space-between;margin:0 12px 12px;text-align:left}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-bN97Pc{background-color:var(--dt-surface,#fff);margin:0}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke{margin:24px 24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke{margin:0}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke-fmcmS{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:1.375rem;font-weight:400;letter-spacing:0;line-height:1.75rem;color:#202124}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-r4nke-fmcmS{background-color:var(--dt-surface,#fff);color:var(--dt-on-surface,#3c4043);font:var(--dt-headline-small-font,400 1.5rem/2rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-headline-small-spacing,0)}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-g7W7Ed{color:#202124;font-family:"Roboto";font-style:normal;font-weight:400;font-size:14px;line-height:20px;letter-spacing:.2px;margin-bottom:22.6px;width:428px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-g7W7Ed{font:var(--dt-body-large-font,400 1rem/1.5rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-large-spacing,0.00625em);margin:24px 0;color:var(--dt-on-surface,#3c4043)}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-c6xFrd{margin-right:22px;margin-left:auto;margin-bottom:18px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;padding:0}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-c6xFrd{margin:0;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;flex-direction:row;width:100%;justify-content:flex-end}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;line-height:20px;border:none;background:#1a73e8;box-sizing:border-box;-moz-border-radius:4px;border-radius:4px;color:#fff;margin:0 12px;min-width:70px;outline:none;padding:8px 24px;text-align:center;cursor:pointer}.ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:14px;line-height:20px;background:#fff;border:1px solid #dadce0;-moz-border-radius:4px;border-radius:4px;box-sizing:border-box;color:#1a73e8;margin:0 12px;min-width:70px;outline:none;padding:8px 24px;text-align:center;cursor:pointer}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe{margin:0 0 0 24px;line-height:20px;-moz-border-radius:100px;border-radius:100px;background:var(--dt-surface,#fff);color:var(--dt-primary,#1a73e8);font:var(--dt-label-large-font,500 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-label-large-spacing,0.0178571429em);border:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe:hover,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe:hover{background:rgba(168,199,250,.08);color:var(--dt-primary,#1a73e8);border:none}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe:focus,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe:focus,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-Rsbfue-LgbsSe:active,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-L7w45e-Rsbfue-LPmGke-Sx9Kwc-IbE0S-LgbsSe:active{background:rgba(168,199,250,.12);color:var(--dt-primary,#1a73e8);border:none;outline:none;-moz-box-shadow:none;box-shadow:none}.ndfHFb-c4YZDc-Wrql6b{background-color:rgba(0,0,0,.6);height:27px;padding:10px 0 10px 0;position:absolute;top:0;width:100%;z-index:3}.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b{background-color:#4d90fe}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b{background-color:rgba(147,147,147,.7);padding:10px 0 10px 0}.ndfHFb-c4YZDc-Wrql6b-hOcTPc{left:20px;position:absolute;white-space:nowrap}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Wrql6b-hOcTPc{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center;position:static}.ndfHFb-c4YZDc-Wrql6b-hOcTPc .ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c{float:right}.ndfHFb-c4YZDc-Wrql6b-LQLjdd{position:absolute;top:0;white-space:nowrap;height:47px}.ndfHFb-c4YZDc-gvZm2b-WAutxc .ndfHFb-c4YZDc-Wrql6b-LQLjdd{background-color:#4d90fe;border-left:1px solid #6aa3ff;border-right:1px solid #6aa3ff}.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-Wrql6b-LQLjdd{border-color:transparent}.ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b{display:inline-block}.ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b{position:absolute;right:16px;top:0;white-space:nowrap}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b{right:0}.ndfHFb-c4YZDc-Wrql6b-N7Eqid{background-color:rgba(0,0,0,.6);display:inline-block;font-size:11px;line-height:28px;margin-right:10px;vertical-align:top}.ndfHFb-c4YZDc-Wrql6b-Bz112c{background-size:contain;display:inline-block;float:left;height:16px;margin-right:12px;position:relative;top:8px;width:16px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-Wrql6b-Bz112c{top:0}.ndfHFb-c4YZDc-Wrql6b-jfdpUb{color:#b3b3b3;display:inline-block}.ndfHFb-c4YZDc-Wrql6b-V1ur5d{color:#fff;font-size:13px;font-weight:normal;line-height:27px}.ndfHFb-c4YZDc-Wrql6b-V1ur5d.ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-qnnXGd{line-height:20px}.ndfHFb-c4YZDc-Wrql6b-V1ur5d-hpYHOb,.ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-hpYHOb{visibility:hidden;position:absolute;height:auto;width:auto}.ndfHFb-c4YZDc-Wrql6b-V1ur5d.ndfHFb-c4YZDc-Iqlsrf-qnnXGd{cursor:pointer}.ndfHFb-c4YZDc-Wrql6b-V1ur5d-hSRGPd:hover{cursor:pointer;text-decoration:underline}.ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d{font-size:11px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b{pointer-events:none;background:linear-gradient(to bottom,rgba(0,0,0,.65) 0%,transparent 100%);height:56px;padding:0 0 16px 0;left:0;right:0;width:auto}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b{height:64px;padding:0;background:transparent}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b.ndfHFb-c4YZDc-Wrql6b-Hyc8Sd{height:64px;padding:0;background:rgba(31,31,31,.85)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-SmKAyb{position:absolute;pointer-events:auto;height:48px;left:0;right:0;padding-top:8px;width:auto}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-SmKAyb{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;justify-content:space-between;align-items:center;padding-top:0;height:64px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b.ndfHFb-c4YZDc-Wrql6b-qbOKL{-moz-box-shadow:0 2px 2px rgba(0,0,0,.6);box-shadow:0 2px 2px rgba(0,0,0,.6);background:#323232;padding:0}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b{background:rgba(0,0,0,.75);height:40px;top:12px;left:auto;padding:0}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b-SmKAyb{height:40px;padding:0;margin:0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{margin-left:8px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-DdWCyb-b0t70b{position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b{top:auto;right:0}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;position:static;align-items:center}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b.ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b-SfQLQb-Woal0c-jcJzye-n1UuX{top:0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-Bz112c{-moz-border-radius:2px;border-radius:2px;margin:3px 11px;width:18px;height:18px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-jfdpUb{letter-spacing:0}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-V1ur5d{font-size:14px;line-height:40px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-V1ur5d{font:var(--dt-title-medium-font,500 1rem/1.5rem "Google Sans"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-title-medium-spacing,0.00625em)}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-V1ur5d.ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-qnnXGd{line-height:30px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-LQLjdd{display:inline-block;position:relative}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-LQLjdd{display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;align-items:center}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-TvD9Pc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{float:left;margin-left:0}.ndfHFb-c4YZDc-hDEnYe{width:100%;height:100%;padding-top:47px;box-sizing:border-box}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-hDEnYe{padding-top:0}.ndfHFb-c4YZDc-i5oIFb:not(.ndfHFb-c4YZDc-e1YmVc) .ndfHFb-c4YZDc-hDEnYe{padding-top:56px}.ndfHFb-c4YZDc-uoC0bf.ndfHFb-c4YZDc-i5oIFb:not(.ndfHFb-c4YZDc-e1YmVc) .ndfHFb-c4YZDc-hDEnYe{padding-top:64px}.ndfHFb-c4YZDc-hDEnYe-SmKAyb{width:100%;height:100%;box-sizing:border-box;padding-bottom:39px}.ndfHFb-c4YZDc-hDEnYe-SmKAyb .ndfHFb-c4YZDc-wvGCSb-gkA7Yd{position:relative;right:initial;top:initial}.ndfHFb-c4YZDc-hDEnYe-AznF2e{width:100%;height:100%;font-size:0;box-sizing:border-box;position:relative}.ndfHFb-c4YZDc-hDEnYe-AznF2e>.ndfHFb-c4YZDc-bN97Pc-u0pjoe-haAclf{position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-hDEnYe-XuHpsb-haAclf{background-color:transparent;z-index:1;overflow:auto;position:absolute;left:0;top:0;right:0;bottom:0}.ndfHFb-c4YZDc-hDEnYe-RwANvf-BvBYQ-haAclf{position:absolute;left:0;bottom:0;overflow-y:hidden}.ndfHFb-c4YZDc-hDEnYe-RwANvf-DKlKme-haAclf{position:absolute;top:0;overflow-x:hidden}.ndfHFb-c4YZDc-hDEnYe-RwANvf-qbOKL-PLDbbf{position:absolute;overflow:hidden}.ndfHFb-c4YZDc-hDEnYe-XuHpsb-qJTHM{position:relative}.ndfHFb-c4YZDc-hDEnYe-Df1ZY-bN97Pc{font-size:11px;opacity:.01;overflow:hidden;position:absolute;width:100%;height:100%;left:0;top:0;z-index:-1;display:block}.ndfHFb-c4YZDc-hDEnYe-fFW7wc{width:100%;z-index:3;background-color:#000;position:absolute;bottom:0;padding-left:46px;box-sizing:border-box;white-space:nowrap;padding-bottom:6px;padding-top:1px}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{font-size:12px;font-weight:normal;padding:0 8px;max-width:200px;overflow:hidden;background-color:#212121;background-image:none;color:#989898;line-height:32px;margin-right:4px;border:none;border-top-right-radius:0;border-top-left-radius:0;border-bottom-right-radius:3px;border-bottom-left-radius:3px;height:inherit;-moz-box-shadow:none;box-shadow:none;text-overflow:ellipsis}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{padding:5px 0 1px 0}.ndfHFb-c4YZDc-hDEnYe-z5C9Gb-Bz112c{background-position:0 -200px;width:24px;height:24px;margin-left:auto;margin-right:auto}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-hDEnYe-z5C9Gb-Bz112c{background-position:0 -2056px}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe{background-color:#4a4a4a;color:white}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-LgbsSe.ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{color:white;cursor:pointer}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob{background-color:#212121;border:none;max-height:200px}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob>.ndfHFb-c4YZDc-j7LFlb{margin:0 20px;padding:0;font-size:12px;color:#989898;height:32px;border:none}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob>.ndfHFb-c4YZDc-j7LFlb>.ndfHFb-c4YZDc-j7LFlb-bN97Pc{max-width:250px;min-width:30px;white-space:nowrap;text-overflow:ellipsis;overflow-x:hidden;line-height:32px;display:inline-block}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob>.ndfHFb-c4YZDc-j7LFlb-sn54Q{color:white;cursor:pointer;background-color:inherit}.ndfHFb-c4YZDc-hDEnYe-fFW7wc-z5C9Gb-xl07Ob>.ndfHFb-c4YZDc-LgbsSe-IwzHHe.ndfHFb-c4YZDc-j7LFlb{background-color:#4a4a4a;color:white}.ndfHFb-c4YZDc-hDEnYe-eFD6re{left:-5000px;position:absolute;top:-5000px}.ndfHFb-c4YZDc-hDEnYe-wvGCSb-gkA7Yd-haAclf .ndfHFb-c4YZDc-wvGCSb-gkA7Yd{left:30px;position:absolute;right:30px;top:0}.ndfHFb-c4YZDc-hDEnYe-wvGCSb-gkA7Yd-haAclf{bottom:39px;overflow:auto;padding-top:8px;position:absolute;left:auto;right:0;top:56px;width:362px}.ndfHFb-c4YZDc-hDEnYe-wvGCSb-bF1uUb{bottom:39px;left:0;overflow:hidden;position:absolute;right:0;top:56px}.ndfHFb-c4YZDc-hDEnYe-jNm5if-Bz112c-awotqb{display:inline-block;margin:0 4px;vertical-align:middle}.ndfHFb-c4YZDc-hDEnYe-jNm5if-NnAfwf-VCkuzd{background:white;-moz-border-radius:2px 2px 0 2px;border-radius:2px 2px 0 2px;color:black;height:16px;min-width:12px;padding:0 4px;position:relative;text-align:center;top:-1px}.ndfHFb-c4YZDc-hDEnYe-jNm5if-NnAfwf{font-family:"Google Sans",Roboto,arial,sans-serif;font-size:10px;position:relative;top:-9px}.ndfHFb-c4YZDc-hDEnYe-jNm5if-Zj4Smb{border-left:4px solid transparent;border-top:4px solid white;height:0;position:absolute;right:0;top:16px;width:0}.ndfHFb-c4YZDc-hDEnYe-wvGCSb-ge6pde-uDEFge{background:#4285f4;left:50%;padding:10px 16px 10px 16px;position:absolute;top:68px;transform:translateX(-50%)}.ndfHFb-c4YZDc-hDEnYe-XuHpsb-hSRGPd-haAclf{-moz-user-select:none}.ndfHFb-c4YZDc-hDEnYe-bN97Pc{position:absolute}.ndfHFb-c4YZDc-fmcmS-RCfa3e{-moz-transition:left .218s ease-out,top .218s ease-out,height .218s ease-out,width .218s ease-out;transition:left .218s ease-out,top .218s ease-out,height .218s ease-out,width .218s ease-out}.ndfHFb-c4YZDc-fmcmS,.ndfHFb-c4YZDc-fmcmS-s2gQvd{bottom:0;position:absolute;top:0;width:100%}.ndfHFb-c4YZDc-fmcmS-haAclf{height:100%;position:absolute;width:100%}.ndfHFb-c4YZDc-fmcmS-s2gQvd{overflow:auto}.ndfHFb-c4YZDc-fmcmS-s2gQvd .ndfHFb-c4YZDc-wvGCSb-gkA7Yd{right:initial}.ndfHFb-c4YZDc-fmcmS-b0t70b{position:absolute}.ndfHFb-c4YZDc-fmcmS-bN97Pc{-moz-user-select:text;background-color:#fff!important;color:#000!important;border:20px solid transparent;font-family:"Courier New",Courier,monospace,arial,sans-serif;font-size:14px;word-wrap:break-word;-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35)}.ndfHFb-c4YZDc-fmcmS-DARUcf{-moz-user-select:text;background-color:#fff!important;color:#000!important;display:block;font-family:"Courier New",Courier,monospace,arial,sans-serif;margin:0;white-space:pre-wrap;word-wrap:break-word}.ndfHFb-c4YZDc-fmcmS-bN97Pc.ndfHFb-c4YZDc-fmcmS-kY93ue,.ndfHFb-c4YZDc-fmcmS-kY93ue .ndfHFb-c4YZDc-fmcmS-DARUcf{-moz-user-select:none;-moz-user-select:none}.ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf{height:100%;position:absolute;width:100%;z-index:1}.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q{position:absolute}.ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c{filter:alpha(opacity=20);opacity:.2;background-color:#28f}.ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd.ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf{filter:alpha(opacity=50);opacity:.5}.ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c{filter:alpha(opacity=40);opacity:.4;background-color:#34a853}.ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-auswjd.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf:not([onclick]):not(:link):not(:visited){background-color:transparent!important}.ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b.ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf{filter:alpha(opacity=.5);opacity:.5}.ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c{filter:alpha(opacity=40);opacity:.4;background-color:#fbbc04}.ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b .ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-auswjd.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-Hl5q5c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-RDNXzf-L6cTce .ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b{display:none}.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q.ndfHFb-c4YZDc-vWsuo-fmcmS-sn54Q-NowJzb{border-bottom:2px solid #fbbc04}.ndfHFb-c4YZDc-JUCs7e{border:3px solid transparent;-moz-border-radius:3px;border-radius:3px;display:inline-block;height:63px;margin:3px 0 3px 3px;outline:none;width:84px}.ndfHFb-c4YZDc-JUCs7e-SmKAyb{display:table-cell;height:inherit;vertical-align:middle;width:inherit}.ndfHFb-c4YZDc-JUCs7e img{display:block;margin:auto}.ndfHFb-c4YZDc-JUCs7e-Bz112c{width:63px;height:63px}.ndfHFb-c4YZDc-JUCs7e-RJLb9c{max-height:63px;max-width:84px}.ndfHFb-c4YZDc-JUCs7e.ndfHFb-c4YZDc-JUCs7e-gk6SMd{border-color:transparent}.ndfHFb-c4YZDc-JUCs7e.ndfHFb-c4YZDc-JUCs7e-ZmdkE,.ndfHFb-c4YZDc-JUCs7e.ndfHFb-c4YZDc-JUCs7e-XpnDCe{border-color:#9c9c9c}.ndfHFb-c4YZDc-q77wGc{position:absolute;left:50%;margin-right:-50%;-moz-transform:translate(-50%);transform:translate(-50%);-moz-border-radius:3px;border-radius:3px;bottom:12px;z-index:3;overflow:hidden}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-q77wGc{-moz-border-radius:100px;border-radius:100px;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex}.ndfHFb-c4YZDc-q77wGc .ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb,.ndfHFb-c4YZDc-q77wGc .ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb{background:rgba(0,0,0,.75)}.ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b .ndfHFb-c4YZDc-LgbsSe.ndfHFb-c4YZDc-C7uZwb-ibnC6b-Btuy5e{-moz-border-radius:25%;border-radius:25%;padding:0}.ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b .ndfHFb-c4YZDc-C7uZwb-ibnC6b-Btuy5e .ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c{transform:scale(0.66667) translateY(-2px)}.ndfHFb-c4YZDc-GSQQnc-LgbsSe,.ndfHFb-c4YZDc-MZArnb-LgbsSe,.ndfHFb-c4YZDc-TvD9Pc-LgbsSe{z-index:1;min-height:24px}.ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{filter:alpha(opacity=87);opacity:0.87;position:relative;margin-left:auto;margin-right:auto}.ndfHFb-c4YZDc-TvD9Pc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-GSQQnc-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-MZArnb-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-DH6Rkf-Bz112c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c,.ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{height:21px;width:21px;margin-top:3px}.ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 0}.ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -1160px}.ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -1280px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-TvD9Pc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -1528px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-MZArnb-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -1712px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-GSQQnc-LgbsSe .ndfHFb-c4YZDc-DH6Rkf-Bz112c{background-position:0 -2304px;height:24px;width:24px;margin:0}.ndfHFb-c4YZDc-i5oIFb.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b .ndfHFb-c4YZDc-GSQQnc-LgbsSe{margin-left:0}.ndfHFb-c4YZDc-tk3N6e-suEOdc.tk3N6e-suEOdc{background-color:#000;border-color:#000;font-family:arial,sans-serif;z-index:1303}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-tk3N6e-suEOdc.tk3N6e-suEOdc{-moz-border-radius:2px;border-radius:2px;font-family:"Google Sans",Roboto,arial,sans-serif}.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-jQ8oHc,.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-jQ8oHc,.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-Ya1KTb .tk3N6e-suEOdc-ez0xG,.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-d6mlqf .tk3N6e-suEOdc-ez0xG{border-color:#000 transparent}.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-jQ8oHc,.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-jQ8oHc,.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-y6n2Me .tk3N6e-suEOdc-ez0xG,.ndfHFb-c4YZDc-tk3N6e-suEOdc .tk3N6e-suEOdc-cX0Lwc .tk3N6e-suEOdc-ez0xG{border-color:transparent #000}.ndfHFb-c4YZDc-neVct-RCfa3e{-moz-transition-property:left,top,width,height;transition-property:left,top,width,height;-moz-transition-duration:.218s;transition-duration:.218s;-moz-transition-timing-function:cubic-bezier(0,0,0.2,1);transition-timing-function:cubic-bezier(0,0,0.2,1)}.ndfHFb-c4YZDc-N4imRe-NMrWyd-RCfa3e{-moz-transition-property:left,right,top,bottom;transition-property:left,right,top,bottom;-moz-transition-duration:.218s;transition-duration:.218s;-moz-transition-timing-function:cubic-bezier(0,0,0.2,1);transition-timing-function:cubic-bezier(0,0,0.2,1)}.ndfHFb-c4YZDc-Wrql6b-zM6fo-GMvhG-b0t70b{display:inline-block}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-Wrql6b-zM6fo-GMvhG-b0t70b{border:1px solid transparent;-moz-border-radius:2px;border-radius:2px;background:rgba(0,0,0,.75);margin:0;white-space:nowrap}.ndfHFb-c4YZDc-zM6fo-GMvhG-Bz112c{background-position:0 -2584px;height:18px;width:18px;margin:2px 4px;position:absolute}.ndfHFb-c4YZDc-zM6fo-GMvhG-fmcmS{line-height:22px;margin:2px 15px 2px 24px;font-size:14px;font-weight:normal}.ndfHFb-c4YZDc-aTv5jf{border:10px solid transparent;position:absolute;z-index:0}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-aTv5jf{border:none}.ndfHFb-c4YZDc-aTv5jf-uquGtd{position:absolute;top:0;left:0;width:100%;height:100%;z-index:1}.ndfHFb-c4YZDc-aTv5jf-AHe6Kc{position:absolute;width:100%;height:100%;top:0;left:0;z-index:1}.ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf{font:13px arial;text-align:center;z-index:2;position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf a{color:#fff!important;text-decoration:underline}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf{color:#1e1e1e}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-aTv5jf-u0pjoe-Ne3sFf a{color:#1e1e1e!important}.ndfHFb-c4YZDc-aTv5jf-bVEB4e{background-color:black;cursor:pointer;position:absolute;top:0;left:0;width:100%;height:100%;z-index:2}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf-NziyQe-Bz112c:not(:link):not(:visited){background-image:url('//ssl.gstatic.com/s2/tt/images/play-overlay.png')!important;background-color:transparent!important;background-repeat:no-repeat;height:77px;width:77px;filter:alpha(opacity=80);opacity:.8}.ndfHFb-c4YZDc-aTv5jf-NziyQe-LgbsSe{z-index:3;filter:alpha(opacity=80);opacity:.8;position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc-aTv5jf-bVEB4e-RJLb9c{height:100%;width:100%}.ndfHFb-c4YZDc:not(.ndfHFb-c4YZDc-e1YmVc) .ndfHFb-c4YZDc-aTv5jf-AHe6Kc{-moz-box-shadow:0px 4px 15px 2px rgba(0,0,0,.35);box-shadow:0px 4px 15px 2px rgba(0,0,0,.35)}.ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde{position:absolute;top:50%;left:50%;margin-right:-50%;-moz-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/v-spinner_dark.gif')!important}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c:not(:link):not(:visited){background-image:none!important}.ndfHFb-c4YZDc .ndfHFb-c4YZDc-aTv5jf .ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS{color:#fff!important}.ndfHFb-c4YZDc-LSZ0mb-fmcmS{margin-left:5px}.ndfHFb-c4YZDc-LSZ0mb-hFsbo{border-left:4px solid transparent;border-right:4px solid transparent;margin-bottom:1px;margin-left:11px;display:inline-block}.ndfHFb-c4YZDc-LSZ0mb-hFsbo-hgHJW{border-top:4px solid rgba(255,255,255,0.87)}.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-LSZ0mb-hFsbo-hgHJW{border-top:4px solid rgba(255,255,255,1)}.ndfHFb-c4YZDc-LSZ0mb-hFsbo-yHKmmc{border-bottom:4px solid rgba(255,255,255,0.87)}.ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-LSZ0mb-hFsbo-yHKmmc{border-bottom:4px solid rgba(255,255,255,1)}.ndfHFb-c4YZDc-kODWGd-xlL3N{height:100%;position:absolute;left:auto;right:10px}.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-LgbsSe{left:-35px;right:auto;position:absolute;top:2px}.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-bMElCd-Bz112c,.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-R6PoUb-Bz112c,.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-ibL1re-Bz112c,.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-c5RTEf-Bz112c{height:28px;width:31px}.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-bMElCd-Bz112c{background-position:0 -2120px}.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-R6PoUb-Bz112c{background-position:0 -2040px}.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-ibL1re-Bz112c{background-position:0 -560px}.ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-c5RTEf-Bz112c{background-position:0 -1400px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-bMElCd-Bz112c{background-position:0 -1408px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-R6PoUb-Bz112c{background-position:0 -3794px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-ibL1re-Bz112c{background-position:0 -2810px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-kODWGd-xlL3N-qPaVXd-r8s4j-c5RTEf-Bz112c{background-position:0 -936px}.ndfHFb-c4YZDc-kODWGd-xlL3N-SxecR{width:40px}.ndfHFb-c4YZDc-kODWGd-xlL3N-SxecR-PFprWc{height:12px;width:12px}.ndfHFb-c4YZDc-deA65-di8rgd-Sx9Kwc{background:#4285f4;-moz-border-radius:2px;border-radius:2px;color:#000;font:normal 13px arial,sans-serif;line-height:20px;position:absolute;width:562px;z-index:1194}.ndfHFb-c4YZDc-deA65-di8rgd-LgbsSe{background:transparent;border:none;color:white;cursor:pointer;float:right;font-size:14px;margin-bottom:auto;margin-left:auto;margin-top:auto;padding:10px 16px;text-decoration:none;text-transform:uppercase}.ndfHFb-c4YZDc-deA65-di8rgd-LgbsSe:hover{outline:white auto 5px}.ndfHFb-c4YZDc-deA65-di8rgd-Sx9Kwc-r4nke-fmcmS,.ndfHFb-c4YZDc-deA65-di8rgd-Sx9Kwc-bN97Pc{float:left;font-size:14px;font-weight:500;padding:10px 32px 10px 16px}.ndfHFb-c4YZDc-nJjxad-nK2kYb,.ndfHFb-c4YZDc-nJjxad-b0t70b{display:inline-block;white-space:nowrap}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-nK2kYb{height:40px}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-nJjxad-b0t70b{margin-left:10px}.ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=87);opacity:0.87;height:21px;width:21px;position:relative;margin-left:auto;margin-right:auto;margin-top:3px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=100);opacity:1;height:24px;width:24px;margin:0}.ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-LgbsSe-OWB6Me .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=47);opacity:0.47}.ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-LgbsSe-ZmdkE .ndfHFb-c4YZDc-Bz112c{filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-nK2kYb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-ZmdkE{background-color:#616161;background-image:none}.ndfHFb-c4YZDc-nJjxad-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -2440px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -776px}.ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe .ndfHFb-c4YZDc-Bz112c{background-position:0 -1360px}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-LgbsSe-IwzHHe .ndfHFb-c4YZDc-Bz112c{background-position:0 -1016px}.ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-nJjxad-ge6pde .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited){background-image:url('//ssl.gstatic.com/docs/common/v-spinner_dark.gif')!important;background-position:0}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-nJjxad-ge6pde .ndfHFb-c4YZDc-Bz112c:not([onclick]):not(:link):not(:visited){background-image:none!important;filter:alpha(opacity=100);opacity:1}.ndfHFb-c4YZDc-vyDMJf-aZ2wEe .ndfHFb-c4YZDc-nJjxad-LgbsSe.ndfHFb-c4YZDc-nJjxad-ge6pde .ndfHFb-aZ2wEe{display:block}.ndfHFb-c4YZDc-nJjxad-SxecR{display:inline-block;height:8px;margin-right:10px;width:100px}.ndfHFb-c4YZDc-nJjxad-SxecR .ndfHFb-c4YZDc-SxecR-skjTt-j4LONd{background-color:#d9d9d9;background-image:-moz-linear-gradient(top,#c3c3c3,#d9d9d9);background-image:linear-gradient(top,#c3c3c3,#d9d9d9);background-color:#d9d9d9!important}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-nJjxad-SxecR .ndfHFb-c4YZDc-SxecR-skjTt-j4LONd{background-color:#fff!important;background-image:none;border-color:transparent!important;-moz-box-shadow:0px 1px 1px 0px rgba(0,0,0,.35);box-shadow:0px 1px 1px 0px rgba(0,0,0,.35)}.ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc{background-color:#151515;background-image:-moz-linear-gradient(top,#000,#303030);background-image:linear-gradient(top,#000,#303030);-moz-box-shadow:0 0 5px 0px #fff;box-shadow:0 0 5px 0px #fff;background-color:#151515!important;-moz-border-radius:6px;border-radius:6px;top:18px;height:10px;width:10px;border:solid 1px #fff}.ndfHFb-c4YZDc-i5oIFb .ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc{top:16px}.ndfHFb-c4YZDc-e1YmVc .ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc{background-color:#58595b!important;background-image:none;height:8px;width:8px;border:solid 2px #fff;margin-left:10px;-moz-box-shadow:0px 1px 1px 0px rgba(0,0,0,.35);box-shadow:0px 1px 1px 0px rgba(0,0,0,.35)}.ndfHFb-c4YZDc-auswjd-gk6SMd .ndfHFb-c4YZDc-SxecR-PFprWc.ndfHFb-c4YZDc-nJjxad-SxecR-PFprWc{background-color:#fff!important;background-image:none;-moz-box-shadow:0px 1px 1px 0px rgba(30,53,69,.9);box-shadow:0px 1px 1px 0px rgba(30,53,69,.9)}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb{display:inline-block;padding:2px;vertical-align:middle}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{-moz-border-radius:1px;border-radius:1px;width:24px;height:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe{-moz-border-radius:100px;border-radius:100px}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe.ndfHFb-c4YZDc-LgbsSe-OWB6Me{filter:alpha(opacity=47);opacity:0.47}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-to915-LgbsSe .ndfHFb-c4YZDc-Bz112c{width:24px;height:24px}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-m9bMae-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -2200px}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-bEDTcc-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -552px}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-hj4D6d-LgbsSe .ndfHFb-c4YZDc-Bz112c{background-position:0 -776px}.ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb .ndfHFb-c4YZDc-nJjxad-hj4D6d-LgbsSe.ndfHFb-c4YZDc-nJjxad-S9gUrf .ndfHFb-c4YZDc-Bz112c{background-position:0 -1016px}.IyROMc-JIbuQc-mJSDk-Bz112c{direction:ltr;text-align:left;overflow:hidden;position:relative;vertical-align:middle}.IyROMc-JIbuQc-mJSDk-RJLb9c:before{content:url(//ssl.gstatic.com/docs/common/shortcut_sprite1.png)}.IyROMc-JIbuQc-mJSDk-RJLb9c{height:95px;position:absolute;width:21px}.IyROMc-JIbuQc-mJSDk-a4fUwd{left:0;top:-63px}.IyROMc-JIbuQc-mJSDk-a4fUwd-HLvlvd{left:0;top:-21px}.IyROMc-JIbuQc-mJSDk-G0jgYd{left:0;top:-42px}.IyROMc-JIbuQc-mJSDk-G0jgYd-HLvlvd{left:0;top:0}.ndfHFb-w37qKe-ppgLk-V68bde{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;vertical-align:middle}.ndfHFb-w37qKe-ppgLk-V68bde-sfGayb-SKd3Ne{margin:auto}.ndfHFb-w37qKe-V68bde{position:absolute;z-index:1002;-moz-box-shadow:rgba(0,0,0,.2) 0 4px 16px;box-shadow:rgba(0,0,0,.2) 0 4px 16px;background-color:#f1f1f1;border:1px solid rgba(0,0,0,.2);color:#6e6e6e;font-size:13px;font-weight:normal;text-align:left;white-space:nowrap}.ndfHFb-w37qKe-V68bde-i5vt6e-L6cTce *:focus{outline:none}.ndfHFb-w37qKe-V68bde-bN97Pc{display:-webkit-box;display:-moz-box;display:-ms-flexbox;display:-webkit-flex;display:flex;padding:10px}.ndfHFb-w37qKe-V68bde-Ne3sFf{overflow:hidden;text-overflow:ellipsis;-webkit-box-orient:vertical;-webkit-line-clamp:6;display:-webkit-box;max-height:90px;margin:auto;max-width:160px;padding-right:10px;word-break:break-word}.ndfHFb-w37qKe-LgbsSe{display:inline-block;margin:auto}.ndfHFb-w37qKe-V68bde-hSRGPd-SKd3Ne{color:#15c;cursor:pointer;padding:0 7px}.ndfHFb-w37qKe-V68bde-TvD9Pc-SKd3Ne{cursor:pointer;height:15px;padding:3px;vertical-align:middle}.ndfHFb-w37qKe-V68bde-hSRGPd-SKd3Ne.ndfHFb-w37qKe-LgbsSe-ZmdkE{text-decoration:underline}.ndfHFb-w37qKe-V68bde-hFsbo{position:absolute;width:20px}.ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe,.ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc{content:"";display:block;height:0;position:absolute;width:0}.ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe{border:10px solid}.ndfHFb-w37qKe-V68bde-hFsbo .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc{border:9px solid}.ndfHFb-w37qKe-V68bde-Ya1KTb{bottom:0}.ndfHFb-w37qKe-V68bde-d6mlqf{top:-10px}.ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe,.ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe{border-color:rgba(0,0,0,.2) transparent;left:0}.ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc,.ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc{border-color:#f1f1f1 transparent;left:1px}.ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe,.ndfHFb-w37qKe-V68bde-Ya1KTb .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc{border-bottom-width:0}.ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-WgXLxe{border-top-width:0}.ndfHFb-w37qKe-V68bde-d6mlqf .ndfHFb-w37qKe-V68bde-Zj4Smb-BuvAkc{border-top-width:0;top:2px}.ndfHFb-w37qKe-Sx9Kwc{-moz-box-shadow:0 4px 16px rgba(0,0,0,.2);box-shadow:0 4px 16px rgba(0,0,0,.2);background:var(--dt-background,#fff);background-clip:padding-box;color:var(--dt-on-surface,#3c4043);font-family:inherit;outline:0;padding:24px;position:absolute;width:560px;z-index:2204}.ndfHFb-w37qKe-Sx9Kwc-xJ5Hnf{background:var(--dt-on-surface,#3c4043);left:0;position:absolute;top:0;z-index:2203}div.ndfHFb-w37qKe-Sx9Kwc-xJ5Hnf{filter:alpha(opacity=50);opacity:.50}.ndfHFb-w37qKe-Sx9Kwc-r4nke{background-color:var(--dt-background,#fff);color:var(--dt-on-surface,#3c4043);cursor:default;font-size:20px;font-weight:normal;line-height:24px}.ndfHFb-w37qKe-Sx9Kwc-r4nke-TvD9Pc{height:11px;margin:24px;opacity:.7;padding:6px;position:absolute;right:0;top:0;width:11px}.ndfHFb-w37qKe-Sx9Kwc-r4nke-TvD9Pc:after{background:url(//ssl.gstatic.com/ui/v1/dialog/close-x.png);content:"";height:11px;position:absolute;width:11px}.ndfHFb-w37qKe-Sx9Kwc-r4nke-TvD9Pc:hover{opacity:1}.ndfHFb-w37qKe-Sx9Kwc-bN97Pc{background-color:var(--dt-background,#fff);font-size:16px;line-height:1.4em;padding-top:24px;padding-bottom:24px;word-wrap:break-word}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd{text-align:right}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe{-moz-border-radius:2px;border-radius:2px;background-color:var(--dt-surface-variant,#f1f3f4);background-image:-moz-linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1);background-image:linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1);border:1px solid #dcdcdc;border:1px solid rgba(0,0,0,.1);color:var(--dt-on-surface,#3c4043);cursor:default;font-family:inherit;font-size:11px;font-weight:bold;height:29px;line-height:27px;margin:0 0 0 16px;min-width:72px;outline:0;padding:0 8px}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe:hover{-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1);background-color:var(--dt-surface-variant,#f1f3f4);background-image:-moz-linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1);background-image:linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1);border:1px solid #c6c6c6;color:var(--dt-on-surface,#3c4043)}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe:active{-moz-box-shadow:0 1px 1px rgba(0,0,0,.1);box-shadow:0 1px 1px rgba(0,0,0,.1);background-color:var(--dt-surface-variant,#f1f3f4);background-image:-moz-linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1);background-image:linear-gradient(top,var(--dt-surface-variant,#f1f3f4),#f1f1f1);border:1px solid #c6c6c6;color:var(--dt-on-surface,#3c4043);-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.1);box-shadow:inset 0 1px 2px rgba(0,0,0,.1)}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe:focus{border:1px solid var(--dt-primary,#1a73e8)}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .ndfHFb-w37qKe-LgbsSe[disabled]{-moz-box-shadow:none;box-shadow:none;background:var(--dt-background,#fff);background-image:none;border:1px solid var(--dt-surface-variant,#f1f3f4);border:1px solid rgba(0,0,0,.5);color:rgba(0,0,0,.26)}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc{background-color:var(--dt-primary,#1a73e8);background-image:-moz-linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8));background-image:linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8));border:1px solid var(--dt-primary,#1a73e8);color:var(--dt-background,#fff)}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:hover{background-color:var(--dt-primary,#1a73e8);background-image:-moz-linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8));background-image:linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8));border:1px solid var(--dt-primary,#1a73e8);color:var(--dt-background,#fff)}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:active{background-color:var(--dt-primary,#1a73e8);background-image:-moz-linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8));background-image:linear-gradient(top,var(--dt-primary,#1a73e8),var(--dt-primary,#1a73e8));border:1px solid var(--dt-primary,#1a73e8);color:var(--dt-background,#fff);-moz-box-shadow:inset 0 1px 2px rgba(0,0,0,.3);box-shadow:inset 0 1px 2px rgba(0,0,0,.3)}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc:focus{-moz-box-shadow:inset 0 0 0 1px #fff;box-shadow:inset 0 0 0 1px #fff;border:1px solid #fff;border:rgba(0,0,0,0) solid 1px;outline:1px solid var(--dt-primary,#1a73e8);outline:rgba(0,0,0,0) 0}.ndfHFb-w37qKe-Sx9Kwc-c6xFrd .VIpgJd-ldDVFe-JIbuQc[disabled]{-moz-box-shadow:none;box-shadow:none;background:var(--dt-primary,#1a73e8);color:var(--dt-background,#fff);filter:alpha(opacity=50);opacity:.5}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-xl07Ob{-moz-box-shadow:none;box-shadow:none;margin-bottom:-24px;padding:0;position:relative;z-index:inherit}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb{color:var(--dt-on-surface,#3c4043);font-size:13px;height:16px;margin:0;opacity:.87;padding:0 0 24px 16px}.ndfHFb-w37qKe-Sx9Kwc-rymPhb-ibnC6b{display:block;overflow:hidden;text-overflow:ellipsis}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-sn54Q{border-left:0;background-color:inherit}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-bN97Pc{margin:0}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-sn54Q .VIpgJd-j7LFlb-bN97Pc,.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-bN97Pc{color:inherit}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-auswjd .VIpgJd-j7LFlb-MPu53c{background:rgba(235,235,235,1)}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-j7LFlb-AHmuwe .VIpgJd-j7LFlb-MPu53c{border-color:var(--dt-primary,#1a73e8)}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-wQNmvb-gk6SMd{background:rgba(255,255,255,0)}.ndfHFb-w37qKe-Sx9Kwc .VIpgJd-wQNmvb-gk6SMd .VIpgJd-j7LFlb-MPu53c::after{-moz-border-radius:50%;border-radius:50%;background:rgba(96,96,96,1);content:"";display:block}.ndfHFb-c4YZDc-SjW3R-ORHb{align-items:center;background:#e8f0fe;color:#202124;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;font-family:"Google Sans",Roboto,arial,sans-serif;height:48px;width:100%}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb{background:#7cacf8;font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-SjW3R-ORHb-haAclf.ndfHFb-c4YZDc-SjW3R-ORHb-L6cTce,.ndfHFb-c4YZDc-SjW3R-ORHb-c6xFrd.ndfHFb-c4YZDc-SjW3R-ORHb-L6cTce,.ndfHFb-c4YZDc-SjW3R-ORHb-L6cTce{display:none}.ndfHFb-c4YZDc-SjW3R-ORHb-c6xFrd{align-items:center;display:-webkit-box;display:-moz-box;display:-webkit-flex;display:-ms-flexbox;display:flex;box-flex:1;flex-grow:1;float:right;justify-content:flex-end}.ndfHFb-c4YZDc-SjW3R-ORHb-Bz112c{background-image:url('//ssl.gstatic.com/docs/common/viewer/v3/v-sprite50.svg');background-position:0 -2722px;height:24px;margin:0 16px;width:24px}.ndfHFb-c4YZDc-SjW3R-ORHb-Ne3sFf{margin-left:16px;font-size:14px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-Ne3sFf{font:var(--dt-body-medium-font,400 .875rem/1.25rem "Roboto"),"Google Sans",Roboto,Arial,sans-serif;letter-spacing:var(--dt-body-medium-spacing,0.0142857143em)}.ndfHFb-c4YZDc-SjW3R-ORHb-IYtByb-LgbsSe-Bz112c{background-position:0 -1160px;height:24px;width:24px}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-IYtByb-LgbsSe-Bz112c{background-position:0 -3570px}.ndfHFb-c4YZDc-SjW3R-ORHb-IYtByb-LgbsSe-sM5MNb{margin:0 16px}.ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe:hover,.ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe:hover{cursor:pointer}.ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe{margin:0 12px;text-align:center;min-width:70px;background:#1a73e8;-moz-border-radius:5px;border-radius:5px;font-size:14px;font-weight:500;padding:7px 0;color:#fff}.ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe:hover{background:#2b7de9}.ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe{margin:0 5px;text-align:center;min-width:70px;color:#1a73e8;font-size:14px;font-weight:500;padding:7px 0}.ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe:hover{background:#f8fbff}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-ssJRIf-LgbsSe:hover,.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-SjW3R-ORHb-K4efff-LgbsSe:hover{background:transparent;color:#202124}.ndfHFb-c4YZDc-zsEIvc-b0t70b{background:white;bottom:0;position:absolute;right:0;top:0;width:320px;z-index:4}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-zsEIvc-b0t70b{background:transparent;-moz-border-radius:24px;border-radius:24px;padding:0 16px 16px 0;box-sizing:border-box;width:344px}.ndfHFb-c4YZDc-zsEIvc-L5Fo6c{border:none;height:100%;width:100%;z-index:4}.ndfHFb-c4YZDc-uoC0bf .ndfHFb-c4YZDc-zsEIvc-L5Fo6c{-moz-border-radius:24px;border-radius:24px}@media only screen and (max-width:500px){.ndfHFb-c4YZDc-zsEIvc-b0t70b{width:100%}}sentinel{}</style></head><body id="yDmH0d" jsmodel="elptZb;PuTOgd" jscontroller="pjICDe" jsaction="rcuQ6b:npT2md; click:FAbpgf; auxclick:FAbpgf;qako4e:.CLIENT;UjQMac:.CLIENT;GvneHb:.CLIENT;c0v8t:.CLIENT;keydown:.CLIENT;keyup:.CLIENT;keypress:.CLIENT;HO6t5b:.CLIENT;mlnRJb:.CLIENT;nHjqDd:.CLIENT" class="tQj5Y ghyPEc IqBfM ecJEib b30Rkd EIlDfe cjGgHb d8Etdd LcUz9d z7HEHd gyaw1d ar1wE UvHKof nTrDbc GAP4ve xSXax AJlUyd CPYzFb V7D6ud fKVgu nk6WKe ndfHFb-c4YZDc-qbOKL-OEVmcd" data-has-header="true" data-no-view="true" style="min-height: 968px;"><script nonce="" aria-hidden="true">window.wiz_progress&&window.wiz_progress();</script><nav jscontroller="Lnriuf" jsaction="tLnfOb:spIfde;qako4e:.CLIENT" class="joJglb" id="kO001e" role="navigation" aria-hidden="true"><div class="QRiHXd"><div class="FXKA9c"><div class="XIpEib QRiHXd"><div class="k43Owe mmOZjd" data-focus-id="JUeBdc"><div><div jscontroller="u6TIZe" jsaction="rcuQ6b:npT2md;JIbuQc:VJ10Y; keydown:I481le;B3adYc:wAhJT" jsmodel="WKE3nf" data-course-states="1" soy-skip="" ssk="5:FHFnz" id="ow4" __is_owner="true"><span data-is-tooltip-wrapper="true"><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc xSP5ic oxacD" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd;" data-idom-class="yHy1rc eT1oJ mN1ivc xSP5ic oxacD" jsname="LgbsSe" aria-label="Menu principal" data-tooltip-enabled="true" data-tooltip-id="tt-i1"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg width="24" height="24" viewBox="0 0 24 24" focusable="false" class=" NMm5M"><path d="M3 18h18v-2H3v2zm0-5h18v-2H3v2zm0-7v2h18V6H3z"></path></svg></span></button><div class="EY8ABd-OWXEXe-TAWMXe" id="tt-i1" role="tooltip" aria-hidden="true">Menu principal</div></span></div></div></div><h1 class="Hwv4mb"><a class="onkcGd OGhwGf" target="_self" href="https://classroom.google.com/c/NTQxMjM1MjY0NzQ5" data-focus-id="/c/NTQxMjM1MjY0NzQ5"><span id="UGb2Qe" class="YVvGBb z3vRcc Pce5Kb">G_MC613B_2023S1</span></a></h1></div></div><div class="R2tE8e QRiHXd VHRSDf "></div><div class="Mtd4hb QRiHXd" soy-skip="" ssk="6:byE9zf"><div class="fB7J9c kWv2Xb QRiHXd"><div style="display: none;"><div jsaction="click:CTftRe" class="XGLVqf oT3cQd" style="display: none;" jsowner="ow724"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD" jsname="KdmTJe" data-tooltip-enabled="true" data-tooltip-override-client-rect="ZAUrGc"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod xSP5ic" aria-hidden="true"><svg enable-background="new 0 0 24 24" focusable="false" height="24" viewBox="0 0 24 24" width="24" class=" NMm5M"><rect fill="none" height="24" width="24"></rect><path d="M7,4L2,9v9c0,1.1,0.9,2,2,2h12c1.1,0,2-0.9,2-2v-4.5l4,4v-11l-4,4V6c0-1.1-0.9-2-2-2H7z M16,18H4v-8l4-4h8V18z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="" target="_blank" aria-label="Participar da videochamada do Meet" data-tooltip-enabled="true" data-tooltip-id="ZAUrGc"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="ZAUrGc">Participar da videochamada do Meet</div></span></div></div><div style="display: none;"><div jsaction="click:CTftRe" class="XGLVqf oT3cQd" style="display: none;" jsowner="ow601"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD" jsname="KdmTJe" data-tooltip-enabled="true" data-tooltip-override-client-rect="ZAUrGc"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod xSP5ic" aria-hidden="true"><svg enable-background="new 0 0 24 24" focusable="false" height="24" viewBox="0 0 24 24" width="24" class=" NMm5M"><rect fill="none" height="24" width="24"></rect><path d="M7,4L2,9v9c0,1.1,0.9,2,2,2h12c1.1,0,2-0.9,2-2v-4.5l4,4v-11l-4,4V6c0-1.1-0.9-2-2-2H7z M16,18H4v-8l4-4h8V18z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="" target="_blank" aria-label="Participar da videochamada do Meet" data-tooltip-enabled="true" data-tooltip-id="ZAUrGc"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="ZAUrGc">Participar da videochamada do Meet</div></span></div></div><div style="display: none;"><div jsaction="rcuQ6b:npT2md;JIbuQc:Ckgp2b(mSMdM);FzgWvd:j697N" class="XGLVqf" jscontroller="RFXpNd" jsowner="ow368"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><span data-is-tooltip-wrapper="true"><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc GR7QId oxacD" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc GR7QId oxacD" jsname="mSMdM" aria-label="Criar ou participar de uma turma" data-tooltip-enabled="true" data-tooltip-id="tt-c6"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 13h-7v7h-2v-7H4v-2h7V4h2v7h7v2z"></path></svg></span></button><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="tt-c6">Criar ou participar de uma turma</div></span></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="true" data-menu-uid="ucc-1"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Adicionar curso&quot;" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="SLuNwd" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Participar da turma</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="svCv4e" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Criar turma</span></li></ul></div></div></div><span data-is-tooltip-wrapper="true"><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc sEZiv TYHMlb oxacD" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc sEZiv TYHMlb oxacD" jsname="mSMdM" aria-label="Participar da turma" data-tooltip-enabled="true" data-tooltip-id="tt-c7"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 13h-7v7h-2v-7H4v-2h7V4h2v7h7v2z"></path></svg></span></button><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="tt-c7">Participar da turma</div></span></div></div><div style="display: none;"><div class="XGLVqf Y5vSD CG2qQ" jsaction="JIbuQc:trigger.FT6KGc" jsowner="ow570"><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD" jsname="dq27Te" aria-label="Configurações da turma" guidedhelpid="courseSettingsGH"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod xSP5ic" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M13.85 22.25h-3.7c-.74 0-1.36-.54-1.45-1.27l-.27-1.89c-.27-.14-.53-.29-.79-.46l-1.8.72c-.7.26-1.47-.03-1.81-.65L2.2 15.53c-.35-.66-.2-1.44.36-1.88l1.53-1.19c-.01-.15-.02-.3-.02-.46 0-.15.01-.31.02-.46l-1.52-1.19c-.59-.45-.74-1.26-.37-1.88l1.85-3.19c.34-.62 1.11-.9 1.79-.63l1.81.73c.26-.17.52-.32.78-.46l.27-1.91c.09-.7.71-1.25 1.44-1.25h3.7c.74 0 1.36.54 1.45 1.27l.27 1.89c.27.14.53.29.79.46l1.8-.72c.71-.26 1.48.03 1.82.65l1.84 3.18c.36.66.2 1.44-.36 1.88l-1.52 1.19c.01.15.02.3.02.46s-.01.31-.02.46l1.52 1.19c.56.45.72 1.23.37 1.86l-1.86 3.22c-.34.62-1.11.9-1.8.63l-1.8-.72c-.26.17-.52.32-.78.46l-.27 1.91c-.1.68-.72 1.22-1.46 1.22zm-3.23-2h2.76l.37-2.55.53-.22c.44-.18.88-.44 1.34-.78l.45-.34 2.38.96 1.38-2.4-2.03-1.58.07-.56c.03-.26.06-.51.06-.78s-.03-.53-.06-.78l-.07-.56 2.03-1.58-1.39-2.4-2.39.96-.45-.35c-.42-.32-.87-.58-1.33-.77l-.52-.22-.37-2.55h-2.76l-.37 2.55-.53.21c-.44.19-.88.44-1.34.79l-.45.33-2.38-.95-1.39 2.39 2.03 1.58-.07.56a7 7 0 0 0-.06.79c0 .26.02.53.06.78l.07.56-2.03 1.58 1.38 2.4 2.39-.96.45.35c.43.33.86.58 1.33.77l.53.22.38 2.55z"></path><circle cx="12" cy="12" r="3.5"></circle></svg></span></button></div></div><div style="display: none;"><div class="XGLVqf Y5vSD CG2qQ" jsaction="JIbuQc:trigger.FT6KGc" jsowner="ow691"><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD" jsname="dq27Te" aria-label="Configurações da turma" guidedhelpid="courseSettingsGH"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod xSP5ic" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M13.85 22.25h-3.7c-.74 0-1.36-.54-1.45-1.27l-.27-1.89c-.27-.14-.53-.29-.79-.46l-1.8.72c-.7.26-1.47-.03-1.81-.65L2.2 15.53c-.35-.66-.2-1.44.36-1.88l1.53-1.19c-.01-.15-.02-.3-.02-.46 0-.15.01-.31.02-.46l-1.52-1.19c-.59-.45-.74-1.26-.37-1.88l1.85-3.19c.34-.62 1.11-.9 1.79-.63l1.81.73c.26-.17.52-.32.78-.46l.27-1.91c.09-.7.71-1.25 1.44-1.25h3.7c.74 0 1.36.54 1.45 1.27l.27 1.89c.27.14.53.29.79.46l1.8-.72c.71-.26 1.48.03 1.82.65l1.84 3.18c.36.66.2 1.44-.36 1.88l-1.52 1.19c.01.15.02.3.02.46s-.01.31-.02.46l1.52 1.19c.56.45.72 1.23.37 1.86l-1.86 3.22c-.34.62-1.11.9-1.8.63l-1.8-.72c-.26.17-.52.32-.78.46l-.27 1.91c-.1.68-.72 1.22-1.46 1.22zm-3.23-2h2.76l.37-2.55.53-.22c.44-.18.88-.44 1.34-.78l.45-.34 2.38.96 1.38-2.4-2.03-1.58.07-.56c.03-.26.06-.51.06-.78s-.03-.53-.06-.78l-.07-.56 2.03-1.58-1.39-2.4-2.39.96-.45-.35c-.42-.32-.87-.58-1.33-.77l-.52-.22-.37-2.55h-2.76l-.37 2.55-.53.21c-.44.19-.88.44-1.34.79l-.45.33-2.38-.95-1.39 2.39 2.03 1.58-.07.56a7 7 0 0 0-.06.79c0 .26.02.53.06.78l.07.56-2.03 1.58 1.38 2.4 2.39-.96.45.35c.43.33.86.58 1.33.77l.53.22.38 2.55z"></path><circle cx="12" cy="12" r="3.5"></circle></svg></span></button></div></div></div><div class="PYWmSe Oe4zIb"><div class="neGRTd"><div class="gb_Fa gb_6d gb_8a gb_Ha" id="gb"><div class="gb_4d gb_6a gb_Sd" ng-non-bindable="" data-ogsr-up=""><div class="gb_Xe"><div class="gb_1c"><div class="gb_N gb_od gb_s gb_Hf" data-ogsr-fb="true" data-ogsr-alt="" id="gbwa"><div class="gb_Ff"><a class="gb_e" aria-label="Google Apps" href="https://www.google.com.br/intl/pt-BR/about/products" aria-expanded="false" role="button" tabindex="0"><svg class="gb_1e" focusable="false" viewBox="0 0 24 24"><path d="M6,8c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2zM12,20c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2zM6,20c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2zM6,14c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2zM12,14c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2zM16,6c0,1.1 0.9,2 2,2s2,-0.9 2,-2 -0.9,-2 -2,-2 -2,0.9 -2,2zM12,8c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2zM18,14c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2zM18,20c1.1,0 2,-0.9 2,-2s-0.9,-2 -2,-2 -2,0.9 -2,2 0.9,2 2,2z"></path></svg></a></div></div></div><div class="gb_b gb_od gb_rg gb_s gb_Hb gb_Hf"><div class="gb_Ff gb_5a gb_rg gb_s"><a class="gb_e gb_1a gb_s" aria-label="Conta do Google: Rafael Andre Alves De Siqueira  
(r243360@dac.unicamp.br)" href="https://accounts.google.com/SignOutOptions?hl=pt-BR&amp;continue=https://classroom.google.com/c/NDQ4MTYxOTM2MzI4" role="button" tabindex="0"><img class="gb_h gbii" src="dec2_to_4_files/unnamed_011.jpg" srcset="dec2_to_4_files/unnamed_011.jpg 1x, dec2_to_4_files/unnamed_013.jpg 2x" alt="" aria-hidden="true" data-noaft=""></a><div class="gb_bb"></div><div class="gb_ab"></div></div></div></div><div style="overflow: hidden; position: absolute; top: 0px; visibility: hidden; width: 328px; z-index: 991; height: 0px; margin-top: 57px; transition: height 0.3s ease-in-out 0s; right: 0px; margin-right: 4px;"><iframe role="presentation" style="height: 100%; width: 100%; visibility: hidden;" scrolling="no" name="app" src="dec2_to_4_files/app.html" frameborder="0"></iframe></div><div style="overflow: hidden; position: absolute; top: 0px; visibility: hidden; width: 400px; z-index: 991; height: 0px; margin-top: 57px; right: 0px; margin-right: 4px;"></div></div></div></div><script nonce="">this.gbar_=this.gbar_||{};(function(_){var window=this;
try{
_.ee=function(a,b,c){if(!a.j)if(c instanceof Array)for(var d of c)_.ee(a,b,d);else{d=(0,_.y)(a.A,a,b);const e=a.s+c;a.s++;b.setAttribute("data-eqid",e);a.B[e]=d;b&&b.addEventListener?b.addEventListener(c,d,!1):b&&b.attachEvent?b.attachEvent("on"+c,d):a.o.log(Error("w`"+b))}};
}catch(e){_._DumpException(e)}
try{
_.fe=function(){if(!_.m.addEventListener||!Object.defineProperty)return!1;var a=!1,b=Object.defineProperty({},"passive",{get:function(){a=!0}});try{_.m.addEventListener("test",()=>{},b),_.m.removeEventListener("test",()=>{},b)}catch(c){}return a}();
}catch(e){_._DumpException(e)}
try{
var ge=document.querySelector(".gb_N .gb_e"),he=document.querySelector("#gb.gb_Rc");ge&&!he&&_.ee(_.Ud,ge,"click");
}catch(e){_._DumpException(e)}
try{
_.wh=function(a){if(a.o)return a.o;for(const b in a.i)if(a.i[b].ta()&&a.i[b].B())return a.i[b];return null};var xh=new class extends _.J{constructor(){var a=_.yc;super();this.B=a;this.o=null;this.j={};this.A={};this.i={};this.s=null}v(a){this.i[a]&&(_.wh(this)&&_.wh(this).K()==a||this.i[a].P(!0))}Ta(a){this.s=a;for(const b in this.i)this.i[b].ta()&&this.i[b].Ta(a)}tc(a){return a in this.i?this.i[a]:null}};_.td("dd",xh);
}catch(e){_._DumpException(e)}
try{
var ij=document.querySelector(".gb_b .gb_e"),jj=document.querySelector("#gb.gb_Rc");ij&&!jj&&_.ee(_.Ud,ij,"click");
}catch(e){_._DumpException(e)}
})(this.gbar_);
// Google Inc.
</script></div></div></div><div class="meR3Qc TeZa2e" jsname="ADG7x"><div class="xHPsid" jsname="njTs3e" role="list"></div></div><div class="WufxEd"></div><div class="QANNMb FJJygb qwLQJ" aria-hidden="false" soy-skip="" ssk="6:bn1bIb"><div class="Olpyd Z3WPhc" aria-live="assertive" aria-atomic="true"></div><div class="tH9B6c Z3WPhc" aria-live="polite" aria-atomic="true"><div style="display: none;"><div class="LhKRUe  " jsowner="ow571" style="display: none;"><span class="dzWTB ">Mural atualizado</span><div class="ar1wZ" jsaction="JIbuQc:aRTGUc"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" aria-label="Mostrar atualizações"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Mostrar</span></button></div></div></div></div><div style="display: none;"><div class="LhKRUe  " jsowner="ow692" style="display: none;"><span class="dzWTB ">Mural atualizado</span><div class="ar1wZ" jsaction="JIbuQc:aRTGUc"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" aria-label="Mostrar atualizações"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Mostrar</span></button></div></div></div></div></div></div><div class="a6pJXc Q6ApZc aTtRxf"><div class="aP3ZPb kRqvHe bFjUmb-Ysl7Fe"><div class="bNpzdf kRqvHe bFjUmb-Wvd9Cc">&nbsp;</div><div class="G1kKid kRqvHe bFjUmb-Wvd9Cc">&nbsp;</div></div></div></nav><div class="FJJygb A2eYae" aria-hidden="true"><div jscontroller="pqmHU" jsaction="rcuQ6b:npT2md;gY980b:B9ntFe" style="display: none" jsmodel="qXV53c" class="Z3WPhc"><div class="LhKRUe  "><span class="dzWTB ">Atualize o navegador para atualizar a página</span><div class="ar1wZ" jsaction="JIbuQc:qrlFte" ssk="9:Atualizar"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd;" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d">Atualizar</span></button></div></div><div class="ar1wZ" jsaction="JIbuQc:IYtByb" ssk="9:Dispensar"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd;" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d">Dispensar</span></button></div></div></div></div><div class="Sslefe Z3WPhc" aria-live="assertive" aria-atomic="true"></div><div class="RmhvCc Z3WPhc" aria-live="polite" aria-atomic="true"></div><div class="w2ifj Z3WPhc" aria-live="polite" aria-atomic="true"><div style="display: none;"><div class="LhKRUe  " style="display: none;"><span class="dzWTB ">Salvando…</span></div></div><div style="display: none;"><div class="LhKRUe  CG2qQ" jsowner="ow593" style="display: none;"><span class="dzWTB ">Você foi convidado a dar aula para esta turma</span><div class="ar1wZ"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me"><div class="VfPpkd-Jh9lGc"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Aceitar</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/invite/accept/NTQxMjI3ODM1NDg1?role=2&amp;continue=%2Fc%2FNTQxMjI3ODM1NDg1&amp;authuser=0" aria-label="Aceitar" data-navigation="server"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div></div></div></div><div style="display: none;"><div class="LhKRUe  D0cJPb" jsowner="ow593"><div class="U51CBd QRiHXd"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20.54 5.23l-1.39-1.68C18.88 3.21 18.47 3 18 3H6c-.47 0-.88.21-1.16.55L3.46 5.23C3.17 5.57 3 6.02 3 6.5V19c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V6.5c0-.48-.17-.93-.46-1.27zM6.24 5h11.52l.83 1H5.42l.82-1zM5 19V8h14v11H5zm11-5.5l-4 4-4-4 1.41-1.41L11 13.67V10h2v3.67l1.59-1.59L16 13.5z"></path></svg></div><span class="dzWTB "><span class="Y5vSD">A turma foi arquivada. Restaure-a para adicionar ou editar informações.</span><span class="nforOe">A turma foi arquivada pelo professor. Não é possível adicionar ou editar informações.</span></span><div class="ar1wZ" jsaction="JIbuQc:E8fGCc"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" aria-label="Restaurar turma arquivada"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Restaurar</span></button></div></div></div></div><div style="display: none;"><div class="LhKRUe  CG2qQ" jsowner="ow714" style="display: none;"><span class="dzWTB ">Você foi convidado a dar aula para esta turma</span><div class="ar1wZ"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me"><div class="VfPpkd-Jh9lGc"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Aceitar</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/invite/accept/NTQxMjM1MjY0NzQ5?role=2&amp;continue=%2Fc%2FNTQxMjM1MjY0NzQ5&amp;authuser=0" aria-label="Aceitar" data-navigation="server"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div></div></div></div><div style="display: none;"><div class="LhKRUe  D0cJPb" jsowner="ow714"><div class="U51CBd QRiHXd"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20.54 5.23l-1.39-1.68C18.88 3.21 18.47 3 18 3H6c-.47 0-.88.21-1.16.55L3.46 5.23C3.17 5.57 3 6.02 3 6.5V19c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V6.5c0-.48-.17-.93-.46-1.27zM6.24 5h11.52l.83 1H5.42l.82-1zM5 19V8h14v11H5zm11-5.5l-4 4-4-4 1.41-1.41L11 13.67V10h2v3.67l1.59-1.59L16 13.5z"></path></svg></div><span class="dzWTB "><span class="Y5vSD">A turma foi arquivada. Restaure-a para adicionar ou editar informações.</span><span class="nforOe">A turma foi arquivada pelo professor. Não é possível adicionar ou editar informações.</span></span><div class="ar1wZ" jsaction="JIbuQc:E8fGCc"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" aria-label="Restaurar turma arquivada"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Restaurar</span></button></div></div></div></div><div style="display: none;"><div class="LhKRUe  CG2qQ" jsowner="ow893" style="display: none;"><span class="dzWTB ">Você foi convidado a dar aula para esta turma</span><div class="ar1wZ"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me"><div class="VfPpkd-Jh9lGc"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Aceitar</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/invite/accept/NTQxMjM1MjY0NzQ5?role=2&amp;continue=%2Fc%2FNTQxMjM1MjY0NzQ5%2Fa%2FNTQzMzAzNDA3NjE3%2Fdetails&amp;authuser=0" aria-label="Aceitar" data-navigation="server"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div></div></div></div><div style="display: none;"><div class="LhKRUe  D0cJPb" jsowner="ow893"><div class="U51CBd QRiHXd"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20.54 5.23l-1.39-1.68C18.88 3.21 18.47 3 18 3H6c-.47 0-.88.21-1.16.55L3.46 5.23C3.17 5.57 3 6.02 3 6.5V19c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V6.5c0-.48-.17-.93-.46-1.27zM6.24 5h11.52l.83 1H5.42l.82-1zM5 19V8h14v11H5zm11-5.5l-4 4-4-4 1.41-1.41L11 13.67V10h2v3.67l1.59-1.59L16 13.5z"></path></svg></div><span class="dzWTB "><span class="Y5vSD">A turma foi arquivada. Restaure-a para adicionar ou editar informações.</span><span class="nforOe">A turma foi arquivada pelo professor. Não é possível adicionar ou editar informações.</span></span><div class="ar1wZ" jsaction="JIbuQc:E8fGCc"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" aria-label="Restaurar turma arquivada"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Restaurar</span></button></div></div></div></div><div><div class="LhKRUe  CG2qQ" jsowner="ow994" style="display: none;"><span class="dzWTB ">Você foi convidado a dar aula para esta turma</span><div class="ar1wZ"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd  U5B3me" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd  U5B3me"><div class="VfPpkd-Jh9lGc"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Aceitar</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/invite/accept/NTQxMjM1MjY0NzQ5?role=2&amp;continue=%2Fc%2FNTQxMjM1MjY0NzQ5%2Fa%2FNTQzMzAzNDAxMzc5%2Fdetails&amp;authuser=0" aria-label="Aceitar" data-navigation="server"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div></div></div></div><div><div class="LhKRUe  D0cJPb" jsowner="ow994"><div class="U51CBd QRiHXd"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20.54 5.23l-1.39-1.68C18.88 3.21 18.47 3 18 3H6c-.47 0-.88.21-1.16.55L3.46 5.23C3.17 5.57 3 6.02 3 6.5V19c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V6.5c0-.48-.17-.93-.46-1.27zM6.24 5h11.52l.83 1H5.42l.82-1zM5 19V8h14v11H5zm11-5.5l-4 4-4-4 1.41-1.41L11 13.67V10h2v3.67l1.59-1.59L16 13.5z"></path></svg></div><span class="dzWTB "><span class="Y5vSD">A turma foi arquivada. Restaure-a para adicionar ou editar informações.</span><span class="nforOe">A turma foi arquivada pelo professor. Não é possível adicionar ou editar informações.</span></span><div class="ar1wZ" jsaction="JIbuQc:E8fGCc"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><button class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 eoooNd Y5vSD U5B3me" aria-label="Restaurar turma arquivada"><div class="VfPpkd-Jh9lGc"></div><div class="VfPpkd-J1Ukfc-LhBDec"></div><div class="VfPpkd-RLmnJb"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Restaurar</span></button></div></div></div></div></div><div class="Ub9MKb Z3WPhc"></div></div><script nonce="" aria-hidden="true">window.wiz_progress&&window.wiz_progress();window.wiz_tick&&window.wiz_tick('BZn5fd');</script><script nonce="" aria-hidden="true">(function(){'use strict';var c=window,d=[];c.aft_counter=d;var e=[],f=0;function _recordIsAboveFold(a){if(!c._isLazyImage(a)&&!a.hasAttribute("data-noaft")&&a.src){var b=(c._isVisible||function(){})(c.document,a);a.setAttribute("data-atf",b);b&&(-1===e.indexOf(a)&&-1===d.indexOf(a)&&d.push(a),a.hasAttribute("data-iml")&&(a=Number(a.getAttribute("data-iml")),a>f&&(f=a)))}}
c.initAft=function(){f=0;e=Array.prototype.slice.call(document.getElementsByTagName("img")).filter(function(a){return!!a.getAttribute("data-iml")});[].forEach.call(document.getElementsByTagName("img"),function(a){try{_recordIsAboveFold(a)}catch(b){throw b.message=a.hasAttribute("data-iid")?b.message+"\nrecordIsAboveFold error for defer inlined image":b.message+("\nrecordIsAboveFold error for img element with <src: "+a.src+">"),b;}});if(0===d.length)c.onaft(f)};}).call(this);
initAft()</script><script id="_ij" nonce="" aria-hidden="true">window.IJ_values = [["112038394563442416565","112038394563442416565","0",false,null,null,true,false], false ,'0','https:\/\/classroom.google.com\/', null ,'boq_apps-edu-classroom-ui_20230313.07_p2','classroom.google.com', 0.0 ,'BR','jDoaUAnrqncRQke8ykU01w','soeYfhSVyVG705UP3dI42A','DEFAULT','', 2023.0 ,'https:\/\/classroom.google.com\/c\/NDQ4MTYxOTM2MzI4', null ,'ltr',[], false , 0.0 ,'\/\/ssl.gstatic.com\/classroom\/favicon.png','https:\/\/accounts.google.com\/AccountChooser?continue\x3dhttps:\/\/classroom.google.com\/c\/NDQ4MTYxOTM2MzI4\x26hl\x3dpt-BR','https:\/\/accounts.google.com\/ServiceLogin?service\x3dclassroom\x26hl\x3dpt-BR\x26authuser\x3d0\x26continue\x3dhttps:\/\/classroom.google.com\/c\/NDQ4MTYxOTM2MzI4','https:\/\/accounts.google.com\/SignOutOptions?continue\x3dhttps:\/\/classroom.google.com\/c\/NDQ4MTYxOTM2MzI4',["https://drive.google.com/picker",null,null,null,null,null,null,null,null,null,null,null,[null,null,"CIvF_fKU_f0CFcdTxAodIq4PLg",1679956297867986,[48475730,48532127,48545168,48548282,45826083,47809549,48642514,47930869,47809351,1787118,47977019,48494755,47893265,47988271,1714246,45814370,47856925,47835375,47860858,1772879,47948077,45754602,45686039,48638933,45775441,1773158,1706538,1729889,48577232,48504704,47807826,48539282,48511759,45771378,1763433,45758671,45774183,48663492,47790498,45735197,48573003,47844885,48410021,49617885,49365716,48475720,48532116,48545154,48548272,45826071,47930858,47809341,48494744,47893254,47988260,47856911,47835361,47948067,45754588,48638923,47807816,48511749,45774169,48663482,47790484,48572993,47844875,49617874,49365706],2],null,null,1000,"",null,null,[null,null,"p",1800000,null,null,null,10000,39000,120000,2,null,100,3100,null,"/punctual/prod/homeroom_prod"],null,null,null,null,null,null,[null,null,"https://gstatic.com/classroom/themes/img_backtoschool.jpg"],null,"r",null,null,null,"",0,null,null,null,null,null,null,null,10,null,null,5,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,10,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,true,null,null,null,null,null,null,null,null,null,null,20,null,null,null,null,null,null,null,null,1000,null,null,"{size}",20,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,"https://calendar.google.com",null,null,null,[100,604800000,2,0.5],null,null,null,null,null,null,null,null,null,null,null,null,null,20,null,null,null,"AIzaSyAewGK8j9KoyT94rEj-weBpysMvzMQzGvk","https://www.googleapis.com/drive/v2internal",null,null,null,null,null,false,null,null,null,true,true,null,null,null,null,null,null,null,null,null,null,null,null,"https://docs.google.com","https://drive.google.com",null,100,null,null,null,null,true,null,"unicamp.br","^video/|^application/(x-flash-video|vnd\\.google-apps\\.video|video)$|^application/vnd\\.google-apps\\.drive-sdk\\.",null,null,null,null,"https://lh3.googleusercontent.com/a/default-user\u003ds72-c-fbw\u003d1",null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,15,null,null,false,null,null,null,null,null,null,false,null,null,null,null,null,null,null,null,null,null,null,null,null,300000,null,null,null,null,null,null,null,10,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,"//ssl.gstatic.com/classroom/favicon.png",null,"30751363934","https://classroom.google.com/",null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,true,null,null,null,4000,1.3,null,null,false,null,[3],null,null,null,null,null,null,null,null,null,null,null,true,null,null,null,null,true,false,null,null,null,null,null,true,null,null,null,null,null,[true,"96485","AIzaSyBqt2sx2fvfwP502G4u_Mu_kRmei_3A2OU",null,false],null,null,null,null,null,false,null,false,null,null,null,null,null,null,null,null,null,200,null,null,null,null,null,null,null,null,null,false,null,null,null,null,null,null,false,null,null,null,null,true,null,null,true,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,true,"BR",null,null,null,null,null,null,["https://workspace.google.com"],null,null,null,null,[false,null,null,null,null,null,null,false,false],null,null,null,null,null,false,null,null,1,null,null,null,false,null,null,null,null,null,null,null,null,null,null,false,null,false,null,1800000,null,null,false,null,null,null,[false,null,[null,null,null,"https://classroom.google.com/ps/create"],true,true],730,null,false,false,false,true,true,false,true,false,false,false,false,false,false,false,false,false,false,false,false], null , false , false , false , false ,'pt','pt-BR',[],'pt_BR','https:\/\/goto2.corp.google.com\/mdtredirect?data_id_filter\x3dclassroom.google.com\x26system_name\x3dapps-edu-classroom-ui', null ,'AD_W2oNDbjunZECTRIvwJkg1TSsp:1679956297868',[["application/vnd.google-apps.document","application/vnd.google-apps.kix"],["application/vnd.google-apps.presentation","application/vnd.google-apps.punch"]], false , null ,'https:\/\/myaccount.google.com\/privacypolicy?hl\x3dpt-BR', false , false ,'https:\/\/myaccount.google.com\/termsofservice?hl\x3dpt-BR','r243360@dac.unicamp.br', true ,'112038394563442416565',]; window.IJ_valuesCb && window.IJ_valuesCb();</script><script id="wiz_jd" nonce="" aria-hidden="true">if (window['_wjdc']) {const wjd = {}; window['_wjdc'](wjd); delete window['_wjdc'];}</script><script id="WIZ-footer" nonce="" aria-hidden="true">window.wiz_progress&&window.wiz_progress(); window.stopScanForCss&&window.stopScanForCss(); ccTick('bl');</script><script nonce="" aria-hidden="true">this.gbar_=this.gbar_||{};(function(_){var window=this;
try{
_.ie=function(a,b){return 0<=_.xb(a,b)};_.je=function(a,b){var c=Array.prototype.slice.call(arguments,1);return function(){var d=c.slice();d.push.apply(d,arguments);return a.apply(this,d)}};_.L=function(a,b){a:if(a=_.E(a,b),null!=a){switch(typeof a){case "string":a=+a;break a;case "number":break a}a=void 0}return a};try{(new self.OffscreenCanvas(0,0)).getContext("2d")}catch(a){};_.ke=function(a,b){this.width=a;this.height=b};_.k=_.ke.prototype;_.k.aspectRatio=function(){return this.width/this.height};_.k.Hb=function(){return!(this.width*this.height)};_.k.ceil=function(){this.width=Math.ceil(this.width);this.height=Math.ceil(this.height);return this};_.k.floor=function(){this.width=Math.floor(this.width);this.height=Math.floor(this.height);return this};_.k.round=function(){this.width=Math.round(this.width);this.height=Math.round(this.height);return this};_.le=function(a,b){return(b||document).getElementsByTagName(String(a))};_.ne=function(a){return _.me(document,a)};_.me=function(a,b){b=String(b);"application/xhtml+xml"===a.contentType&&(b=b.toLowerCase());return a.createElement(b)};_.oe=function(a){for(var b;b=a.firstChild;)a.removeChild(b)};_.pe=function(a){return 9==a.nodeType?a:a.ownerDocument||a.document};
}catch(e){_._DumpException(e)}
try{
var He;_.Fe=function(a,b){if(void 0!==a.i||void 0!==a.j)throw Error("B");a.j=b;_.Ld(a)};_.Ge=class extends _.I{constructor(a){super(a)}};He=0;_.Ke=function(a){return Object.prototype.hasOwnProperty.call(a,_.nb)&&a[_.nb]||(a[_.nb]=++He)};_.Le=function(a){return _.vd(_.rd.i(),a)};
}catch(e){_._DumpException(e)}
try{
_.nj=function(a,b,c){a.rel=c;-1!=c.toLowerCase().indexOf("stylesheet")?(a.href=_.Ic(b),(b=_.id(a.ownerDocument&&a.ownerDocument.defaultView))&&a.setAttribute("nonce",b)):a.href=b instanceof _.Gc?_.Ic(b):b instanceof _.Kc?_.Lc(b):_.Lc(_.Tc(b))};
}catch(e){_._DumpException(e)}
try{
_.oj=function(a){const b=_.Ec();a=b?b.createScriptURL(a):a;return new _.Gc(a,_.Fc)};/*

 SPDX-License-Identifier: Apache-2.0
*/
var pj;try{new URL("s://g"),pj=!0}catch(a){pj=!1}_.qj=pj;
}catch(e){_._DumpException(e)}
try{
_.rj=function(a){var b;let c;const d=null==(c=(b=(a.ownerDocument&&a.ownerDocument.defaultView||window).document).querySelector)?void 0:c.call(b,"script[nonce]");(b=d?d.nonce||d.getAttribute("nonce")||"":"")&&a.setAttribute("nonce",b)};
}catch(e){_._DumpException(e)}
try{
var sj=function(a,b,c){_.Td.log(46,{att:a,max:b,url:c})},uj=function(a,b,c){_.Td.log(47,{att:a,max:b,url:c});a<b?tj(a+1,b):_.yc.log(Error("Y`"+a+"`"+b),{url:c})},tj=function(a,b){if(vj){const d=_.ne("SCRIPT");d.async=!0;d.type="text/javascript";d.charset="UTF-8";var c=d;c.src=_.Hc(vj);_.rj(c);d.onload=_.je(sj,a,b,d.src);d.onerror=_.je(uj,a,b,d.src);_.Td.log(45,{att:a,max:b,url:d.src});_.le("HEAD")[0].appendChild(d)}},wj=class extends _.I{constructor(a){super(a)}};var xj=_.G(_.Od,wj,17)||new wj,yj,vj=(yj=_.G(xj,_.sc,1))?_.oj(_.E(yj,4)||""):null,zj,Aj=(zj=_.G(xj,_.sc,2))?_.oj(_.E(zj,4)||""):null,Bj=function(){tj(1,2);if(Aj){const a=_.ne("LINK");a.setAttribute("type","text/css");_.nj(a,Aj,"stylesheet");let b=_.id();b&&a.setAttribute("nonce",b);_.le("HEAD")[0].appendChild(a)}};(function(){const a=_.Pd();if(_.F(a,18))Bj();else{const b=_.L(a,19)||0;window.addEventListener("load",()=>{window.setTimeout(Bj,b)})}})();
}catch(e){_._DumpException(e)}
})(this.gbar_);
// Google Inc.
</script><div ng-non-bindable="" aria-hidden="true"></div><div jscontroller="mdfgKd" jsaction="rcuQ6b:rcuQ6b;qako4e:rcuQ6b;aWRkAb:pwuS5c;qFdNBb:Pb2hxc;" jsmodel="Var0bb" role="contentinfo" class="dkQQje" guidedhelpid="helpMenuGH" style="" aria-hidden="true"><div role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;;keydown:I481le;" jsshadow="" jsname="LgbsSe" aria-label="Ajuda e comentários" aria-disabled="false" tabindex="0" data-tooltip="Ajuda e comentários" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-menu-corner="bottom-start" data-anchor-corner="top-start" data-tooltip-position="right" data-tooltip-vertical-offset="0" data-tooltip-horizontal-offset="-12"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg width="24" height="24" viewBox="0 0 24 24" focusable="false" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span></span></div></div><div class="gb_Qd" ng-non-bindable="" aria-hidden="true">Google Apps</div><div class="gb_k" ng-non-bindable="" aria-hidden="true"><div class="gb_zc"><div>Conta do Google</div><div class="gb_yb">Rafael Andre Alves De Siqueira</div><div>r243360@dac.unicamp.br</div></div></div><script nonce="" aria-hidden="true">window['HqyC7b'] = window.performance && performance.timing.navigationStart + performance.now();</script><div jsaction="rcuQ6b:npT2md; click:okAHKe(GGAcbc); keydown:I481le;ZldWJd:FNFY6c;zsYKuc:YdzvGf" class="vhK44c dgqqXe" jscontroller="pWaBX" jsowner="ow4" aria-hidden="true"><div class="AxPfNe" jsname="GGAcbc"></div><div class="ETRkCe" jsname="haAclf"><div class="Du1LZe" jscontroller="nW2QJc" jsaction="rcuQ6b:rcuQ6b; click:YdzvGf(ibnC6b); keydown:I481le;lHU8dd:rcuQ6b;qako4e:rcuQ6b;NBlzmd:bQDp8;FZ977b:rcuQ6b"><div class="OX4Vcb" role="menu"><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/h" aria-label="Turmas " role="menuitem" href="https://classroom.google.com/h"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="JDxyrc xSP5ic"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 3L4 9v12h16V9l-8-6zm6 16h-3v-6H9v6H6v-9l6-4.5 6 4.5v9z"></path></svg></div><div class="kXvNXe"><div class="asQXV YVvGBb">Turmas</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/calendar/this-week/course/all" aria-label="Agenda " role="menuitem" href="https://classroom.google.com/calendar/this-week/course/all"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="JDxyrc xSP5ic"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 4h-1V2h-2v2H8V2H6v2H5c-1.11 0-1.99.9-1.99 2L3 20a2 2 0 0 0 2 2h14c1.1 0 2-.9 2-2V6c0-1.1-.9-2-2-2zm0 16H5V9h14v11z"></path></svg></div><div class="kXvNXe"><div class="asQXV YVvGBb">Agenda</div></div></a><li role="separator" class="VfPpkd-rymPhb-clz4Ic e6pQl yCa5be"></li><div role="section" aria-label="Inscrito"><div class="pkktJb iLjzDc YVvGBb">Inscrito</div><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/a/not-turned-in/all" aria-label="Pendentes " role="menuitem" href="https://classroom.google.com/a/not-turned-in/all"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="JDxyrc xSP5ic"><svg enable-background="new 0 0 24 24" focusable="false" height="24" viewBox="0 0 24 24" width="24" class=" NMm5M"><g><rect fill="none" height="24" width="24"></rect></g><g><g><path d="M20,3H4C2.9,3,2,3.9,2,5v14c0,1.1,0.9,2,2,2h16c1.1,0,2-0.9,2-2V5 C22,3.9,21.1,3,20,3z M20,19H4V5h16V19z" fill-rule="evenodd"></path><polygon fill-rule="evenodd" points="19.41,10.42 17.99,9 14.82,12.17 13.41,10.75 12,12.16 14.82,15"></polygon><rect fill-rule="evenodd" height="2" width="5" x="5" y="7"></rect><rect fill-rule="evenodd" height="2" width="5" x="5" y="11"></rect><rect fill-rule="evenodd" height="2" width="5" x="5" y="15"></rect></g></g></svg></div><div class="kXvNXe"><div class="asQXV YVvGBb">Pendentes</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NTQzMjI4NzkxNzU0" aria-label="MC322AB - Programação Orientada a Objetos " role="menuitem" data-id="543228791754" href="https://classroom.google.com/c/NTQzMjI4NzkxNzU0"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  Ag4wUb"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">M</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">MC322AB - Programação Orientada a Objetos</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NTQxMjI3ODM1NDg1" aria-label="G_CE304C_2023S1 " role="menuitem" data-id="541227835485" href="https://classroom.google.com/c/NTQxMjI3ODM1NDg1"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  ee1HBc"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_CE304C_2023S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NTQxMjM0OTIyNTcw" aria-label="G_EE533A_2023S1 " role="menuitem" data-id="541234922570" href="https://classroom.google.com/c/NTQxMjM0OTIyNTcw"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  ee1HBc"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_EE533A_2023S1</div></div></a><a class="Xi8cpb qs41qe" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NTQxMjM1MjY0NzQ5" aria-label="G_MC613B_2023S1 " role="menuitem" data-id="541235264749" href="https://classroom.google.com/c/NTQxMjM1MjY0NzQ5"><div class="LlcfK bFjUmb-Ysl7Fe"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  UvHKof"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_MC613B_2023S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NTI2MjIyODY5MzE1" aria-label="G_CE838A_2022S2 " role="menuitem" data-id="526222869315" href="https://classroom.google.com/c/NTI2MjIyODY5MzE1"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  ee1HBc"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_CE838A_2022S2</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NTM3ODgzMzY5MTQ1" aria-label="G_CE738A_2022S2 " role="menuitem" data-id="537883369145" href="https://classroom.google.com/c/NTM3ODgzMzY5MTQ1"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  UvHKof"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_CE738A_2022S2</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NDQ4MTYxOTM2MzI4" aria-label="G_MC202A+B+C_2022S1 " role="menuitem" data-id="448161936328" href="https://classroom.google.com/c/NDQ4MTYxOTM2MzI4"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  ee1HBc"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_MC202A+B+C_2022S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NDU4MDk2MTg3NDMy" aria-label="G_EE400A_2022S1 " role="menuitem" data-id="458096187432" href="https://classroom.google.com/c/NDU4MDk2MTg3NDMy"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  WFUiUb"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_EE400A_2022S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/NDU4MTAyNTE1ODIy" aria-label="G_F 315A_2022S1 " role="menuitem" data-id="458102515822" href="https://classroom.google.com/c/NDU4MTAyNTE1ODIy"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  UvHKof"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_F 315A_2022S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/Mzc0MzkxMzI3NzQ1" aria-label="G_MC504A_2021S2 " role="menuitem" data-id="374391327745" href="https://classroom.google.com/c/Mzc0MzkxMzI3NzQ1"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  S3aLQd"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_MC504A_2021S2</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/MjYzMDkxODIwMzc4" aria-label="G_EA513A_2021S1 " role="menuitem" data-id="263091820378" href="https://classroom.google.com/c/MjYzMDkxODIwMzc4"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  S3aLQd"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_EA513A_2021S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/MjYzMTMxNjk1NDI5" aria-label="G_F 315A_2021S1 " role="menuitem" data-id="263131695429" href="https://classroom.google.com/c/MjYzMTMxNjk1NDI5"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  ee1HBc"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_F 315A_2021S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/MjY0Nzk4MTgxMTc3" aria-label="G_MS211D_2021S1 " role="menuitem" data-id="264798181177" href="https://classroom.google.com/c/MjY0Nzk4MTgxMTc3"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  ee1HBc"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">G</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">G_MS211D_2021S1</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/c/MjY0NzU0NTEzNTY0" aria-label="HZ291B_2021S1 " role="menuitem" data-id="264754513564" href="https://classroom.google.com/c/MjY0NzU0NTEzNTY0"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="yXVLvd"><div class="CNpREd  S3aLQd"><div aria-hidden="true" class="vUBwW TGnLfc A6dC2c UISY8d-Tvm9db bFjUmb-Tvm9db">H</div></div></div><div class="kXvNXe"><div class="asQXV YVvGBb">HZ291B_2021S1</div></div></a></div><li role="separator" class="VfPpkd-rymPhb-clz4Ic e6pQl yCa5be"></li><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/h/archived" aria-label="Turmas arquivadas " role="menuitem" href="https://classroom.google.com/h/archived"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="JDxyrc xSP5ic"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20.54 5.23l-1.39-1.68C18.88 3.21 18.47 3 18 3H6c-.47 0-.88.21-1.16.55L3.46 5.23C3.17 5.57 3 6.02 3 6.5V19c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V6.5c0-.48-.17-.93-.46-1.27zM6.24 5h11.52l.83 1H5.42l.82-1zM5 19V8h14v11H5zm11-5.5l-4 4-4-4 1.41-1.41L11 13.67V10h2v3.67l1.59-1.59L16 13.5z"></path></svg></div><div class="kXvNXe"><div class="asQXV YVvGBb">Turmas arquivadas</div></div></a><a class="Xi8cpb" jsname="ibnC6b" tabindex="-1" data-focus-id="/s" aria-label="Configurações " role="menuitem" href="https://classroom.google.com/s"><div class="LlcfK"><div class="p1KYTc"></div></div><div class="JDxyrc xSP5ic"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M13.85 22.25h-3.7c-.74 0-1.36-.54-1.45-1.27l-.27-1.89c-.27-.14-.53-.29-.79-.46l-1.8.72c-.7.26-1.47-.03-1.81-.65L2.2 15.53c-.35-.66-.2-1.44.36-1.88l1.53-1.19c-.01-.15-.02-.3-.02-.46 0-.15.01-.31.02-.46l-1.52-1.19c-.59-.45-.74-1.26-.37-1.88l1.85-3.19c.34-.62 1.11-.9 1.79-.63l1.81.73c.26-.17.52-.32.78-.46l.27-1.91c.09-.7.71-1.25 1.44-1.25h3.7c.74 0 1.36.54 1.45 1.27l.27 1.89c.27.14.53.29.79.46l1.8-.72c.71-.26 1.48.03 1.82.65l1.84 3.18c.36.66.2 1.44-.36 1.88l-1.52 1.19c.01.15.02.3.02.46s-.01.31-.02.46l1.52 1.19c.56.45.72 1.23.37 1.86l-1.86 3.22c-.34.62-1.11.9-1.8.63l-1.8-.72c-.26.17-.52.32-.78.46l-.27 1.91c-.1.68-.72 1.22-1.46 1.22zm-3.23-2h2.76l.37-2.55.53-.22c.44-.18.88-.44 1.34-.78l.45-.34 2.38.96 1.38-2.4-2.03-1.58.07-.56c.03-.26.06-.51.06-.78s-.03-.53-.06-.78l-.07-.56 2.03-1.58-1.39-2.4-2.39.96-.45-.35c-.42-.32-.87-.58-1.33-.77l-.52-.22-.37-2.55h-2.76l-.37 2.55-.53.21c-.44.19-.88.44-1.34.79l-.45.33-2.38-.95-1.39 2.39 2.03 1.58-.07.56a7 7 0 0 0-.06.79c0 .26.02.53.06.78l.07.56-2.03 1.58 1.38 2.4 2.39-.96.45.35c.43.33.86.58 1.33.77l.53.22.38 2.55z"></path><circle cx="12" cy="12" r="3.5"></circle></svg></div><div class="kXvNXe"><div class="asQXV YVvGBb">Configurações</div></div></a></div></div></div></div><div id="goog-lr-70" style="position: absolute; top: -1000px; height: 1px; overflow: hidden;" aria-live="polite" aria-atomic="true" aria-hidden="true">LAB03</div><iframe id="hfcr" style="display: none;" src="dec2_to_4_files/RotateCookiesPage.html" aria-hidden="true"></iframe><c-wiz c-wiz="" jsrenderer="g1e71c" class="SSPGKf fXYYpf oCHqfe JwkDRc BIIBbc" jsdata="deferred-c5" data-p="%.@.[1,3],[1,2]]" jscontroller="gQQbc" jsaction="rcuQ6b:rcuQ6b;HO6t5b:PlQWd;gHPzkc:jsAJsc;QmtCl:.CLIENT;qVp5ue:.CLIENT;AE9bOd:.CLIENT;mlnRJb:.CLIENT;lHU8dd:.CLIENT" data-node-index="0;0" jsmodel="hc6Ubd PuTOgd;IaLzN;U9kKWe;WKE3nf;aMcbid;lkzLle;elptZb;" data-ogpc="" data-view-id="ucc-0" data-primary-model="true" data-course-states="1,3" data-course-ready-states="1,2" data-include-abusive-courses="true" style="visibility: hidden; opacity: 0; position: fixed; inset: 0px 0px -1417px; display: none;" aria-busy="true" data-savescroll="0" aria-hidden="true"><div jsname="a9kxte" class="T4LgNb "><div jsname="qJTHM" class="kFwPee"><div class="xgkURe mhCMAe"></div><div class="xgkURe ECPFEb"></div><div jsaction="rcuQ6b:rcuQ6b" jscontroller="FRimSc"></div><div jsaction="rcuQ6b:rcuQ6b;JIbuQc:hskLsf(ZUkOIc); click:RByGDd(XTYNyb)" role="region" jscontroller="V8Zje" aria-label="Banner informativo" aria-hidden="true"></div><div class="bg6sud" jscontroller="AthZQc" jsaction="rcuQ6b:rcuQ6b;lHU8dd:rcuQ6b" jsmodel="WKE3nf" data-course-states="1"><div class="xtiq3"><div jsaction="rcuQ6b:rcuQ6b;FZ977b:rcuQ6b" jscontroller="s3KsTb"></div><div jsaction="rcuQ6b:rcuQ6b;FZ977b:rcuQ6b" jscontroller="I2RHf"></div></div><div class="xtiq3 N33kHb"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 pOf0gc UJYYgf n42Gr VfPpkd-ksKsZd-mWPk3d" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 pOf0gc UJYYgf n42Gr"><div class="VfPpkd-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg enable-background="new 0 0 24 24" focusable="false" height="18" viewBox="0 0 24 24" width="18" class=" NMm5M"><g><rect fill="none" height="24" width="24"></rect></g><g><g><path d="M20,3H4C2.9,3,2,3.9,2,5v14c0,1.1,0.9,2,2,2h16c1.1,0,2-0.9,2-2V5 C22,3.9,21.1,3,20,3z M20,19H4V5h16V19z" fill-rule="evenodd"></path><polygon fill-rule="evenodd" points="19.41,10.42 17.99,9 14.82,12.17 13.41,10.75 12,12.16 14.82,15"></polygon><rect fill-rule="evenodd" height="2" width="5" x="5" y="7"></rect><rect fill-rule="evenodd" height="2" width="5" x="5" y="11"></rect><rect fill-rule="evenodd" height="2" width="5" x="5" y="15"></rect></g></g></svg></span><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Pendentes</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/a/not-turned-in/all" aria-label="Pendentes"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc nQaZq LgeCif xSP5ic" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc nQaZq LgeCif xSP5ic" data-tooltip-enabled="true" data-tooltip-override-client-rect="yfL0u"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><svg enable-background="new 0 0 24 24" focusable="false" height="24" viewBox="0 0 24 24" width="24" class=" NMm5M"><g><rect fill="none" height="24" width="24"></rect></g><g><g><path d="M20,3H4C2.9,3,2,3.9,2,5v14c0,1.1,0.9,2,2,2h16c1.1,0,2-0.9,2-2V5 C22,3.9,21.1,3,20,3z M20,19H4V5h16V19z" fill-rule="evenodd"></path><polygon fill-rule="evenodd" points="19.41,10.42 17.99,9 14.82,12.17 13.41,10.75 12,12.16 14.82,15"></polygon><rect fill-rule="evenodd" height="2" width="5" x="5" y="7"></rect><rect fill-rule="evenodd" height="2" width="5" x="5" y="11"></rect><rect fill-rule="evenodd" height="2" width="5" x="5" y="15"></rect></g></g></svg><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/a/not-turned-in/all" aria-label="Pendentes" data-tooltip-enabled="true" data-tooltip-id="yfL0u"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="yfL0u">Pendentes</div></span><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 pOf0gc UJYYgf n42Gr VfPpkd-ksKsZd-mWPk3d" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 pOf0gc UJYYgf n42Gr"><div class="VfPpkd-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="18" height="18" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 4h-1V2h-2v2H8V2H6v2H5c-1.11 0-1.99.9-1.99 2L3 20a2 2 0 0 0 2 2h14c1.1 0 2-.9 2-2V6c0-1.1-.9-2-2-2zm0 16H5V9h14v11z"></path></svg></span><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Agenda</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/calendar/this-week/course/all" aria-label="Agenda"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc nQaZq LgeCif xSP5ic" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc nQaZq LgeCif xSP5ic" data-tooltip-enabled="true" data-tooltip-override-client-rect="g7hDSd"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 4h-1V2h-2v2H8V2H6v2H5c-1.11 0-1.99.9-1.99 2L3 20a2 2 0 0 0 2 2h14c1.1 0 2-.9 2-2V6c0-1.1-.9-2-2-2zm0 16H5V9h14v11z"></path></svg><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/calendar/this-week/course/all" aria-label="Agenda" data-tooltip-enabled="true" data-tooltip-id="g7hDSd"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="g7hDSd">Agenda</div></span></div></div><div jscontroller="aXmj4" jsaction="rcuQ6b:rcuQ6b;IKbv3d:rcuQ6b;wJx4ze:rcuQ6b;Vgg7gc:yMMCof;iZo7Zb:u2HSyd;yyauTb:.CLIENT;ymHzQd:.CLIENT" jsmodel="I8BbUd;QJeGre;RH7Ihb;qwZZpc"><div jscontroller="CJc2td" jsname="CCJ0ld" data-drag-list-group-key="1" data-drag-direction-left-right="true"><ol jsname="bN97Pc" class="JwPp0e"><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="543228791754" data-user-id="30751363934" data-course-id="543228791754"><div class="Tc9hUd CNpREd Ag4wUb"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_reachout.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQzMjI4NzkxNzU0"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NTQzMjI4NzkxNzU0" data-focus-id="/c/NTQzMjI4NzkxNzU0"><div class="YVvGBb z3vRcc-ZoZQ1">MC322AB - Programação Orientada a Objetos</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQzMjI4NzkxNzU0"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-2"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Esther Luna Colombini</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_009.jpg" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb543228791754" data-focus-id="PMg5Xd-543228791754"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NTQzMjI4NzkxNzU0/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;MC322AB - Programação Orientada a Objetos&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb543228791754" jsaction=""></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb543228791754">Abrir seu trabalho para "MC322AB - Programação Orientada a Objetos"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe543228791754"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/1lm3WuryI4KekSdm1xw4lpraJoPoH91TU0HrASGwHjd95R6Gh7j4isNOtyjx3xaRGvOvOtMIn?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;MC322AB - Programação Orientada a Objetos&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe543228791754" jsaction=""></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe543228791754">Abrir a pasta de "MC322AB - Programação Orientada a Objetos" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="541227835485" data-user-id="30751363934" data-course-id="541227835485"><div class="Tc9hUd CNpREd ee1HBc"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_graduation.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQxMjI3ODM1NDg1"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NTQxMjI3ODM1NDg1" data-focus-id="/c/NTQxMjI3ODM1NDg1"><div class="YVvGBb z3vRcc-ZoZQ1">G_CE304C_2023S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQxMjI3ODM1NDg1"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-3"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Luis Renato Vedovato</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_005.png" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb541227835485" data-focus-id="PMg5Xd-541227835485"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NTQxMjI3ODM1NDg1/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_CE304C_2023S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb541227835485" jsaction=""></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb541227835485">Abrir seu trabalho para "G_CE304C_2023S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe541227835485"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/1lTJUPba_b9tuPoLMjaepVmRq27gpj0fuYeFu5mWDj4F158Nj1BQjwQl2IcXTFLIJJJchWweZ?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_CE304C_2023S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe541227835485"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe541227835485">Abrir a pasta de "G_CE304C_2023S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="541234922570" data-user-id="30751363934" data-course-id="541234922570"><div class="Tc9hUd CNpREd ee1HBc"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_backtoschool.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQxMjM0OTIyNTcw"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NTQxMjM0OTIyNTcw" data-focus-id="/c/NTQxMjM0OTIyNTcw"><div class="YVvGBb z3vRcc-ZoZQ1">G_EE533A_2023S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQxMjM0OTIyNTcw"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-4"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Pedro Xavier de Oliveira</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_002.jpg" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb541234922570" data-focus-id="PMg5Xd-541234922570"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NTQxMjM0OTIyNTcw/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_EE533A_2023S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb541234922570" jsaction=""></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb541234922570">Abrir seu trabalho para "G_EE533A_2023S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe541234922570"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/1BVxXaIvmxftFAYd_NCfYylhMrvrxTESd5tPeTSJIRHYwXC4l67PuGPQp-BIkzB2lpwTYhbjw?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_EE533A_2023S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe541234922570"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe541234922570">Abrir a pasta de "G_EE533A_2023S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="541235264749" data-user-id="30751363934" data-course-id="541235264749"><div class="Tc9hUd CNpREd UvHKof"><div class="OjOEXb" style="background-image: url(&quot;https://lh3.googleusercontent.com/hr_crs_themes/AOy-etcoLWshMMuOyuEPi6my1-CGqcB9Xu_JtMHnnqanhyxe6G4JBb0c4t4iCXmTVmGELBHr5m1J3yZjKSy54B4J-1t-DexpdAV-6W6fpizt1pTinEKhdc5iWqk=s1280&quot;);"></div><div class="ZizeYd bFjUmb-Tvm9db"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQxMjM1MjY0NzQ5"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NTQxMjM1MjY0NzQ5" data-focus-id="/c/NTQxMjM1MjY0NzQ5"><div class="YVvGBb z3vRcc-ZoZQ1">G_MC613B_2023S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTQxMjM1MjY0NzQ5"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-5"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Ricardo Pannain</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_008.jpg" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb541235264749" data-focus-id="PMg5Xd-541235264749"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NTQxMjM1MjY0NzQ5/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_MC613B_2023S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb541235264749" jsaction=""></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb541235264749">Abrir seu trabalho para "G_MC613B_2023S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe541235264749"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/1xc8yZQHDxLusvVvUGlJb563t31KQR-7XjVOljaU2xfvClpG3w-NuPqXT3GIDZKO3LeXhTYCt?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_MC613B_2023S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe541235264749"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe541235264749">Abrir a pasta de "G_MC613B_2023S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="526222869315" data-user-id="30751363934" data-course-id="526222869315"><div class="Tc9hUd CNpREd ee1HBc"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_backtoschool.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTI2MjIyODY5MzE1"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NTI2MjIyODY5MzE1" data-focus-id="/c/NTI2MjIyODY5MzE1"><div class="YVvGBb z3vRcc-ZoZQ1">G_CE838A_2022S2</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTI2MjIyODY5MzE1"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-6"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Marcelo Pereira da Cunha</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_005.jpg" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb526222869315" data-focus-id="PMg5Xd-526222869315"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NTI2MjIyODY5MzE1/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_CE838A_2022S2&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb526222869315"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb526222869315">Abrir seu trabalho para "G_CE838A_2022S2"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe526222869315"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/1l9ZgDX1JWad338Q_yqF8wllcZURR10a-zP4FBQPtqpYkRLVcD6Kc1cX-ISTlj_CLkBixhI3B?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_CE838A_2022S2&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe526222869315"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe526222869315">Abrir a pasta de "G_CE838A_2022S2" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="537883369145" data-user-id="30751363934" data-course-id="537883369145"><div class="Tc9hUd CNpREd UvHKof"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_read.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTM3ODgzMzY5MTQ1"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NTM3ODgzMzY5MTQ1" data-focus-id="/c/NTM3ODgzMzY5MTQ1"><div class="YVvGBb z3vRcc-ZoZQ1">G_CE738A_2022S2</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NTM3ODgzMzY5MTQ1"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-7"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Mauricio Aguiar Serra</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_005.png" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb537883369145" data-focus-id="PMg5Xd-537883369145"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NTM3ODgzMzY5MTQ1/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_CE738A_2022S2&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb537883369145"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb537883369145">Abrir seu trabalho para "G_CE738A_2022S2"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe537883369145"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/18VTbZ2QecASSykuBqf5MVK1Qac6S91L4cwB8eAPqy8k99j2oU4nf1R4NmW8cgBqtSdKXlGxA?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_CE738A_2022S2&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe537883369145"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe537883369145">Abrir a pasta de "G_CE738A_2022S2" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="448161936328" data-user-id="30751363934" data-course-id="448161936328"><div class="Tc9hUd CNpREd ee1HBc"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_graduation.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NDQ4MTYxOTM2MzI4"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NDQ4MTYxOTM2MzI4" data-focus-id="/c/NDQ4MTYxOTM2MzI4"><div class="YVvGBb z3vRcc-ZoZQ1">G_MC202A+B+C_2022S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NDQ4MTYxOTM2MzI4"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-8"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">ORLANDO LEE</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_005.png" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb448161936328" data-focus-id="PMg5Xd-448161936328"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NDQ4MTYxOTM2MzI4/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_MC202A+B+C_2022S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb448161936328"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb448161936328">Abrir seu trabalho para "G_MC202A+B+C_2022S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe448161936328"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/12v5aOOWUCLRVqRQixZjsu-EdVbtA1ydyJu0GQ2GZUl1g6NlXEhzSYXowNiR9MVXB7mi7qyEQ?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_MC202A+B+C_2022S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe448161936328"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe448161936328">Abrir a pasta de "G_MC202A+B+C_2022S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="458096187432" data-user-id="30751363934" data-course-id="458096187432"><div class="Tc9hUd CNpREd WFUiUb"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_bookclub.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NDU4MDk2MTg3NDMy"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NDU4MDk2MTg3NDMy" data-focus-id="/c/NDU4MDk2MTg3NDMy"><div class="YVvGBb z3vRcc-ZoZQ1">G_EE400A_2022S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NDU4MDk2MTg3NDMy"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-9"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">João Bosco Ribeiro do Val</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_005.png" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb458096187432" data-focus-id="PMg5Xd-458096187432"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NDU4MDk2MTg3NDMy/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_EE400A_2022S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb458096187432"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb458096187432">Abrir seu trabalho para "G_EE400A_2022S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe458096187432"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/1x9QcXIyT9LIkbtWHOSneIE_Qv21kcbefpkl6gufXciUQsVjsySwHOAgJE7sk63rmaI55gyZY?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_EE400A_2022S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe458096187432"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe458096187432">Abrir a pasta de "G_EE400A_2022S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="458102515822" data-user-id="30751363934" data-course-id="458102515822"><div class="Tc9hUd CNpREd UvHKof"><div class="OjOEXb" style="background-image: url(&quot;https://lh3.googleusercontent.com/hr_crs_themes/AOy-etdyloexyH3r1hNZDagQFoF7GGoGgmSQKm_VvcXjAj13pyNh4IfhfxVKSD_saWl3PHQdLIqRG9mLw97LnXBYIWDPufiMaoxz1Febcf4hrS1ll8qC_Br1BIU=s1280&quot;);"></div><div class="ZizeYd bFjUmb-Tvm9db"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NDU4MTAyNTE1ODIy"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/NDU4MTAyNTE1ODIy" data-focus-id="/c/NDU4MTAyNTE1ODIy"><div class="YVvGBb z3vRcc-ZoZQ1">G_F 315A_2022S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/NDU4MTAyNTE1ODIy"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-10"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Antonio Vidiella Barranco</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_004.jpg" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb458102515822" data-focus-id="PMg5Xd-458102515822"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/NDU4MTAyNTE1ODIy/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_F 315A_2022S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb458102515822"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb458102515822">Abrir seu trabalho para "G_F 315A_2022S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe458102515822"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/1YNt8oV2mzo2pBpB9sA7GWR4EUrjidgQ-WMSjPbIpjBqHiJjDTAxByBaLoaqvY6G3pWcvi9Mh?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_F 315A_2022S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe458102515822"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe458102515822">Abrir a pasta de "G_F 315A_2022S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="374391327745" data-user-id="30751363934" data-course-id="374391327745"><div class="Tc9hUd CNpREd S3aLQd"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_reachout.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/Mzc0MzkxMzI3NzQ1"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/Mzc0MzkxMzI3NzQ1" data-focus-id="/c/Mzc0MzkxMzI3NzQ1"><div class="YVvGBb z3vRcc-ZoZQ1">G_MC504A_2021S2</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/Mzc0MzkxMzI3NzQ1"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-11"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Arthur Catto</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_002.png" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb374391327745" data-focus-id="PMg5Xd-374391327745"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/Mzc0MzkxMzI3NzQ1/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_MC504A_2021S2&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb374391327745"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb374391327745">Abrir seu trabalho para "G_MC504A_2021S2"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe374391327745"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/17QQRa8U2KXgwW4EApM_D84kCly6lSKXlacyWSra0_cbPnRYYNMoqMiyVefpP34nbpcMyrfVq?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_MC504A_2021S2&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe374391327745"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe374391327745">Abrir a pasta de "G_MC504A_2021S2" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="263091820378" data-user-id="30751363934" data-course-id="263091820378"><div class="Tc9hUd CNpREd S3aLQd"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_reachout.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjYzMDkxODIwMzc4"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/MjYzMDkxODIwMzc4" data-focus-id="/c/MjYzMDkxODIwMzc4"><div class="YVvGBb z3vRcc-ZoZQ1">G_EA513A_2021S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjYzMDkxODIwMzc4"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-12"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Akebo Yamakami</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_005.png" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb263091820378" data-focus-id="PMg5Xd-263091820378"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/MjYzMDkxODIwMzc4/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_EA513A_2021S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb263091820378"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb263091820378">Abrir seu trabalho para "G_EA513A_2021S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe263091820378"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/0B3XmWde0ZxzNflFwdjdQTkl6X19pc2pKam5ZYkE5MzNDQ3FjTkpmTGphU2t6aUItVnd5bDQ?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_EA513A_2021S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe263091820378"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe263091820378">Abrir a pasta de "G_EA513A_2021S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="263131695429" data-user-id="30751363934" data-course-id="263131695429"><div class="Tc9hUd CNpREd ee1HBc"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_graduation.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjYzMTMxNjk1NDI5"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/MjYzMTMxNjk1NDI5" data-focus-id="/c/MjYzMTMxNjk1NDI5"><div class="YVvGBb z3vRcc-ZoZQ1">G_F 315A_2021S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjYzMTMxNjk1NDI5"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-13"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Lázaro Aurélio Padilha</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed.jpg" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb263131695429" data-focus-id="PMg5Xd-263131695429"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/MjYzMTMxNjk1NDI5/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_F 315A_2021S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb263131695429"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb263131695429">Abrir seu trabalho para "G_F 315A_2021S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe263131695429"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/0B3XmWde0ZxzNfkowN1dyYzIwS0RkUEtYZWpWYVdEZnNzX2lHYUliVk12N2JvSmlOOHg4NlU?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_F 315A_2021S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe263131695429"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe263131695429">Abrir a pasta de "G_F 315A_2021S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="264798181177" data-user-id="30751363934" data-course-id="264798181177"><div class="Tc9hUd CNpREd ee1HBc"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_graduation.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjY0Nzk4MTgxMTc3"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/MjY0Nzk4MTgxMTc3" data-focus-id="/c/MjY0Nzk4MTgxMTc3"><div class="YVvGBb z3vRcc-ZoZQ1">G_MS211D_2021S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjY0Nzk4MTgxMTc3"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-14"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Peter Sussner</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_005.png" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb264798181177" data-focus-id="PMg5Xd-264798181177"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/MjY0Nzk4MTgxMTc3/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;G_MS211D_2021S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb264798181177"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb264798181177">Abrir seu trabalho para "G_MS211D_2021S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe264798181177"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/0B3XmWde0ZxzNfm8zaWNBSkI1WVVEZ1BSTlRvUjZLV2ExZ3NSRTBDSU5JZGFMei1ldktNdGs?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;G_MS211D_2021S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe264798181177"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe264798181177">Abrir a pasta de "G_MS211D_2021S1" no Google Drive</div></span></div></div></li><li jsmodel="hCpsVc bYzLLb AKq4rd" class="gHz6xd Aopndd rZXyy" data-draggable-item-id="264754513564" data-user-id="30751363934" data-course-id="264754513564"><div class="Tc9hUd CNpREd S3aLQd"><div class="O7utsb bFjUmb-Tvm9db"></div><div class="OjOEXb Gf8MK" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_reachout.jpg&quot;);"></div><div class="R4EiSb"><a class="onkcGd ZmqAt Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjY0NzU0NTEzNTY0"></a><h2 class="prWPdf"><a class="onkcGd eDfb1d YVvGBb Vx8Sxd" target="_self" href="https://classroom.google.com/c/MjY0NzU0NTEzNTY0" data-focus-id="/c/MjY0NzU0NTEzNTY0"><div class="YVvGBb z3vRcc-ZoZQ1">HZ291B_2021S1</div><div class="YVvGBb"></div></a><a class="onkcGd Nmpzvc Vx8Sxd" target="_self" aria-hidden="true" tabindex="-1" href="https://classroom.google.com/c/MjY0NzU0NTEzNTY0"> </a><div jscontroller="gZb3ib" jsaction="FzgWvd:j697N" data-guided-help-id="courseCardActionMenuGH"><div jsaction="JIbuQc:aj0Jcf(WjL7X); keydown:uYT2Vb(WjL7X);iFFCZc:oNPcuf;Rld2oe:li9Srb" jsshadow="" class="VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd" jscontroller="wg1P6b" jsname="pzCKEc"><div jsname="WjL7X" jsslot=""><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc oxacD JRosVd" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc oxacD JRosVd" aria-label="Opções da turma"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></button></div><div jsname="U0exHf" jsslot=""> <div class="VfPpkd-xl07Ob-XxIAqe VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL VfPpkd-xl07Ob q6oraf P77izf" jscontroller="ywOR5c" jsaction="keydown:I481le;JIbuQc:j697N(rymPhb);XVaHYd:c9v4Fb(rymPhb);Oyo5M:b5fzT(rymPhb);DimkCe:TQSy7b(rymPhb);m0LGSd:fAWgXe(rymPhb);WAiFGd:kVJJuc(rymPhb)" data-is-hoisted="false" data-should-flip-corner-horizontally="false" data-menu-uid="ucc-15"><ul class="VfPpkd-StrnGf-rymPhb DMZ54e" jsname="rymPhb" jscontroller="PHUIyb" jsaction="mouseleave:JywGue; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; keydown:I481le" role="menu" tabindex="-1" aria-label="Menu &quot;Opções&quot; da turma" data-disable-idom="true"><span aria-hidden="true" class="VfPpkd-BFbNVe-bF1uUb NZp2ef"></span><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="QEskHf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Mover</span></li><li class=" VfPpkd-StrnGf-rymPhb-ibnC6b" jsaction="click:o6ZaF;keydown:RDtNu; keyup:JdS61c; focusin:MeMJlc; focusout:bkTmIf;mousedown:teoBgf; mouseup:NZPHBc; mouseenter:SKyDAe; mouseleave:xq3APb; touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8; change:uOgbud" role="menuitem" jsname="ytavkf" tabindex="-1" data-menu-item-skip-restore-focus="true"><span class="VfPpkd-StrnGf-rymPhb-pZXsl"></span><span jsname="K4r5Ff" class="VfPpkd-StrnGf-rymPhb-b9t22c">Cancelar inscrição</span></li></ul></div></div></div></div></h2><div class="QRiHXd"><div class="Vx8Sxd YVvGBb jJIbcc">Pedro Peixoto Ferreira</div><div class="lJv9ke"></div></div></div></div><div class="TQYOZc"><img class="PNzAWd" aria-hidden="true" src="dec2_to_4_files/unnamed_010.jpg" data-atf="false"><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div></div></div><div class="SZ0kZe"><div data-guided-help-id="courseCardStudentProfileGH"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" data-tooltip-enabled="true" data-tooltip-override-client-rect="zxtDBb264754513564" data-focus-id="PMg5Xd-264754513564"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1s-2.4.84-2.82 2H5c-1.1 0-2 .9-2 2v14c0 1.1.9 2 2 2h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7.55 0c.14-.15.33-.25.55-.25s.41.1.55.25c.12.13.2.31.2.5 0 .41-.34.75-.75.75s-.75-.34-.75-.75c0-.19.08-.37.2-.5zM19 5v10.79C16.52 14.37 13.23 14 12 14s-4.52.37-7 1.79V5h14zM5 19v-.77C6.74 16.66 10.32 16 12 16s5.26.66 7 2.23V19H5z"></path><path d="M12 13c1.94 0 3.5-1.56 3.5-3.5S13.94 6 12 6 8.5 7.56 8.5 9.5 10.06 13 12 13zm0-5c.83 0 1.5.67 1.5 1.5S12.83 11 12 11s-1.5-.67-1.5-1.5S11.17 8 12 8z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://classroom.google.com/c/MjY0NzU0NTEzNTY0/sp/MzA3NTEzNjM5MzRa/all" aria-label="Abrir seu trabalho para &quot;HZ291B_2021S1&quot;" data-tooltip-enabled="true" data-tooltip-id="zxtDBb264754513564"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="zxtDBb264754513564">Abrir seu trabalho para "HZ291B_2021S1"</div></span></div><div jscontroller="N8q7Ze" jsaction="rcuQ6b:rcuQ6b;RwVyRc:rcuQ6b"><span data-is-tooltip-wrapper="true"><div class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc eaBpBc" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc eaBpBc" data-tooltip-enabled="true" data-tooltip-override-client-rect="pUkKFe264754513564"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><span class="VfPpkd-kBDsod" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M20 6h-8l-2-2H4c-1.1 0-1.99.9-1.99 2L2 18c0 1.1.9 2 2 2h16c1.1 0 2-.9 2-2V8c0-1.1-.9-2-2-2zm0 12H4V8h16v10z"></path></svg></span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6" href="https://drive.google.com/drive/folders/0B3XmWde0ZxzNfmRVVFdyYVZMOFFSUVdsSTdxU0xCaXliMGhIZ3k3S094aFdDM3ByZVZtdW8?authuser=0" target="_blank" aria-label="Abrir a pasta de &quot;HZ291B_2021S1&quot; no Google Drive" data-tooltip-enabled="true" data-tooltip-id="pUkKFe264754513564"></a><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div></div><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="pUkKFe264754513564">Abrir a pasta de "HZ291B_2021S1" no Google Drive</div></span></div></div></li></ol></div></div><div jscontroller="cs6ocd" jsaction="rcuQ6b:npT2md;FttMgb:Qp7hp;qFdNBb:Pb2hxc;Cvbxce:N6n54b;mlnRJb:p5Uonb" style="display: none;" data-wait-for="aXmj4"></div><div jscontroller="ISr1Vb" jsaction="qFdNBb:Pb2hxc;Cvbxce:ysXIce;lHU8dd:pcE7Z;rcuQ6b:npT2md;FZ977b:pcE7Z" jsmodel="WKE3nf" data-course-states="2" id="ow368" __is_owner="true"></div></div></div><c-data id="c5"></c-data><view-header style="display: none;"><title>Turmas</title></view-header></c-wiz><div id="goog-lr-370" style="position: absolute; top: -1000px; height: 1px; overflow: hidden;" aria-live="assertive" aria-atomic="true" aria-hidden="true"></div><c-wiz c-wiz="" jsrenderer="BZn5fd" class="SSPGKf fXYYpf JwkDRc oCHqfe BIIBbc" jsdata="deferred-c8" data-p="%.@.&quot;NTQxMjI3ODM1NDg1&quot;]" jscontroller="gQQbc" jsaction="rcuQ6b:rcuQ6b;HO6t5b:PlQWd;gHPzkc:jsAJsc;QmtCl:.CLIENT;qVp5ue:.CLIENT;AE9bOd:.CLIENT;mlnRJb:.CLIENT;uwjiC:.CLIENT" data-node-index="0;0" jsmodel="hc6Ubd PuTOgd;IaLzN;U9kKWe;bYzLLb;lkzLle;" data-ogpc="" data-view-id="ucc-16" data-include-user-lists="true" data-course-states="1" style="visibility: hidden; opacity: 0; position: fixed; inset: 0px 0px -772px; display: none;" aria-busy="true" data-savescroll="0" aria-hidden="true"><div jsname="a9kxte" class="T4LgNb "><div jsname="qJTHM" class="kFwPee"><div class="xgkURe mhCMAe"></div><div class="xgkURe ECPFEb"></div><div jsaction="rcuQ6b:rcuQ6b" jscontroller="FRimSc"></div><div jsaction="rcuQ6b:rcuQ6b;JIbuQc:hskLsf(ZUkOIc); click:RByGDd(XTYNyb)" role="region" jscontroller="V8Zje" aria-label="Banner informativo" aria-hidden="true"></div><div class="dbEQNc"><div jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:Fmspve(Q7N4Oc);KAD0te:O99HCf" jscontroller="KHqDY" jsmodel="hb3e8b" class="v9TZ3c bFjUmb-Tvm9db"><div class="qyN25"><div class="PFLqgc PagUde" style="background-image: url(&quot;https://gstatic.com/classroom/themes/img_graduation.jpg&quot;);"><div class="VVnuU ra2NV ee1HBc"></div></div><div class="T4tcpe PagUde"><h1 class="tNGpbb YrFhrf-ZoZQ1 YVvGBb">G_CE304C_2023S1</h1><div class="qFmcrc z3vRcc-ZoZQ1 YVvGBb"></div></div></div></div><div class="M7zXZd"><aside role="complementary" class="DXLeqd"><div class="CG2qQ dsW6Nd"><div jscontroller="UqV0cb" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b"><div jscontroller="RO1Frf" jsaction="rcuQ6b:rcuQ6b;rKHbQd:r2JIKb;HGIkz:VlevBc;uwjiC:rcuQ6b;JIbuQc:RYcsse(BIFOEb)" class="d4Fe0d LBlAUc NA2Gt" style="display: none;" id="ow601" __is_owner="true"><div class="NGVAIb QRiHXd"><img src="dec2_to_4_files/logo_meet_2020q4_color_1x_web_48dp.png" alt="" aria-hidden="true" class="RponAc" data-atf="false"><span class="asQXV">Meet</span><div class="fPqOAb"></div><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb oxacD" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" aria-label="Opções do link do Meet" aria-disabled="false" tabindex="0" aria-haspopup="true" aria-expanded="false" data-alignright="true"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span><div jsname="xl07Ob" style="display: none;" aria-hidden="true"><div role="menu" tabindex="0" class="JPdR6b hVNH5c" jscontroller="uY3Nvd" jsaction="IpSVtb:TvD9Pc;fEN2Ze:xzS4ub;frq95c:LNeFm;cFpp9e:J9oOtd; click:H8nU8b; mouseup:H8nU8b; keydown:I481le; keypress:Kr2w4b; blur:O22p3e; focus:H8nU8b"><div class="XvhY1d" jsaction="mousedown:p8EH2c; touchstart:p8EH2c"><div class="JAPqpe K0NPx"></div></div></div></div></div></div></div></div><div jscontroller="UqV0cb" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b"></div><div class="d4Fe0d LBlAUc "><div class="WMQb5e" jsmodel="hCpsVc"><h2 class="EZrbnd sxa9Pc">Próximas atividades</h2><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div><div class="CHJgKd"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 uBUej n42Gr" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 uBUej n42Gr"><div class="VfPpkd-Jh9lGc"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Ver tudo</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/a/not-turned-in/NTQxMjI3ODM1NDg1" aria-label="Ver todas as atividades"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div></div></div></div></div></div></aside><main class="Sgw65b kdAl3b" jsmodel="uJydvc;I8BbUd;UvJ3Mb;" tabindex="-1" role="main"><div jsmodel="NYdJ9b" data-include-stream-item-materials="false" data-stream-item-types="3" data-list-type="5" data-active-filter="1" data-load-all-pages="true"><div jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;oquPK:rcuQ6b;o2F6Cf:if3DMb" jscontroller="s2wDwf"></div></div><section guidedhelpid="streamContentGH" role="section" jsmodel="NYdJ9b" data-include-stream-item-materials="false" data-list-type="3" data-active-filter="2" data-load-all-pages="false"><div jsaction="rcuQ6b:BU4fHd;HO6t5b:BU4fHd;oquPK:E3Ktff;uwjiC:E3Ktff,rcuQ6b;wJx4ze:rcuQ6b;gbLJWc:ZLWxKf;JIbuQc:fyRA7e(idVoDf);gY980b:B9ntFe" jscontroller="yidvwe" id="ow571" __is_owner="true"><div jscontroller="fJcHcd" class="zOtZye LBlAUc GWZ7yf nmFHZb" jsaction="rcuQ6b:rcuQ6b;peFp2d:Fck3Oe;QAK2O:huHkmc;M6YzAd:Bv9PPc"><div class="zTrXGf "><div class="qk0lee QRiHXd VBEdtc-Wvd9Cc" jsaction="click:Fck3Oe" tabindex="0" role="button" guidedhelpid="courseInlineCreatorGH"><div class="U2zcIf"><div jscontroller="tF6Lzd" jsaction="rcuQ6b:rcuQ6b;FZ977b:rcuQ6b"><img class="tkmmwb" jsname="xJzy8c" aria-hidden="true" src="dec2_to_4_files/unnamed_007.jpg" data-atf="false" width="40px" height="40px"></div></div><div class="K6Ovqd">Escreva um aviso para sua turma</div></div><div class="Y5vSD fidHdf" jsaction="JIbuQc:pJN26"><span data-is-tooltip-wrapper="true"><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" jsname="JC5QVe" aria-label="Reutilizar postagem" data-tooltip-enabled="true" data-tooltip-id="tt-c11" guidedhelpid="courseReuseGH"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod xSP5ic" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 5H4v6h2V7h13M5 19h15v-6h-2v4H5"></path><path d="M16.29 10.71l-1.41-1.42L18.17 6l-3.29-3.29 1.41-1.42L21 6zm-8.58 12L3 18l4.71-4.71 1.41 1.42L5.83 18l3.29 3.29z"></path></svg></span></button><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="tt-c11">Reutilizar postagem</div></span></div></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543876597714" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;Direito e Moral&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "Direito e Moral"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Luis Renato Vedovato postou uma nova atividade: Direito e Moral</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 23 de mar.</span><span aria-hidden="true">23 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543876597714" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 26 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 26 dias.</div></div><div><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543876597714" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543876597714"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543876597714"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543876641332" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;Início da Personalidade Jurídica&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "Início da Personalidade Jurídica"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Luis Renato Vedovato postou uma nova atividade: Início da Personalidade Jurídica</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 23 de mar.</span><span aria-hidden="true">23 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543876641332" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 26 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 26 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543876641332" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543876641332"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543876641332"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543542460825" class="qhnNic LBlAUc Aopndd TIunU"><div class="n4xnA"><div class="JZicYb QRiHXd"><img class="tnyRnb tkmmwb" aria-hidden="true" src="dec2_to_4_files/unnamed_003.png" data-atf="false"><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Aviso: "Equality within Our Lifetimes: How Laws…"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Luis Renato Vedovato</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 14 de mar.</span><span aria-hidden="true">14 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543542460825" data-tooltip=" Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 17 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 17 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="false" data-show-bump="true" data-stream-item-id="543542460825" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Oções de aviso"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div><div class="n8F6Jd"><div class="pco8Kc obylVb j70YMc"><span>Equality within Our Lifetimes: How Laws and Policies Can Close – or Widen – Gender Gaps in Economies Worldwide<br>se puderem baixar esse texto, será ótimo. debate sobre a igualdade.&nbsp;<br><a target="_blank" href="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide">https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide</a></span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;wuANJc:.CLIENT;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel="PTCFbe hGbFme BrMJ0e" data-stream-item-id="543542460825" data-is-edit-mode="false" data-filter="0" data-material-parent-id="PTCFbe" data-include-stream-item-materials="true"><div jsname="UYewLd" class="AgzMgb rhFKgc" style=""><div jsaction="rcuQ6b:rcuQ6b;KtPeHe:rcuQ6b;wuANJc:rcuQ6b" jscontroller="TPuMf" data-parent-id="PTCFbe" jsname="C2Qrw"></div><div class="MlZb9c d3aYgd " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;IKzbTb:Yo3LPb;wuANJc:.CLIENT" jsname="C2Qrw" data-parent-id="PTCFbe" data-mode="7" data-copies-only="false" data-show-originality-analyses="false" data-forms-only="false" data-read-only="false"><div class="luto0c" data-dom-id="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide-0-1-4-https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide-Events &amp; Launches - WORLD Policy Analysis Center-$$-false-false-false-false-$-$-https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide"><a class="VkhHKd e7EEH nQaZq" target="_blank" aria-label="Anexo: link para https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" jsaction="LWntbc" href="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" data-focus-id="eTkQDe-https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" data-attachment-id="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" jsname="HzV7m" data-dom-id="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide-0-1-4-https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide-Events &amp; Launches - WORLD Policy Analysis Center-$$-false-false-false-false-$-$-https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide"><div class="DAnlhb bFjUmb-Wvd9Cc"></div><div class="gM4mlb bFjUmb-Wvd9Cc"></div><div class="rzTfPe xSP5ic "><span class="DPvwYc" aria-hidden="true"></span></div><div class="lIHx8b YVvGBb asQXV ">Events &amp; Launches - WORLD Policy Analysis Center</div></a><div class="pOf0gc QRiHXd Aopndd M4LFnf" jsname="XgfUnd" data-attachment-id="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" jsaction="JIbuQc:Rsbfue(Rsbfue);"><a class="vwNuXe JkIgWb QRiHXd MymH0d maXJsd" target="_blank" aria-label="Anexo: link para https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" jsaction="LWntbc" href="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" title="Events &amp; Launches - WORLD Policy Analysis Center" data-focus-id="hSRGPd-auswjd-https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide-https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide" data-attachment-id="https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide"><div class="bxp7vf bHOAdb Niache"><img jsname="q4uQmd" jsaction="error:dyBsCf" class=" " src="dec2_to_4_files/unnamed_012.jpg" aria-hidden="true" role="presentation" data-mime-type="" data-atf="false"></div><div class="MM30Lb"><div class="A6dC2c QDKOcc VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">Events &amp; Launches - WORLD Policy Analysis Center</div><div class="cSyPgb WInaFd QRiHXd"><div class="QRiHXd"><div class="kRYv9b YVvGBb">https://www.worldpolicycenter.org/events-launches/equality-within-our-lifetimes-how-laws-and-policies-can-close-or-widen-gender-gaps-in-economies-worldwide</div></div></div></div></a><div class="ZgfM9 QRiHXd"></div></div></div></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="MlZb9c d3aYgd " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="7" data-material-parent-id="PTCFbe"></div></div></div><div jsname="QkPyvd" class="" style="display: none;"></div></div></div></div><div role="region" jsname="EQPzXb" class="s2g3Xd "><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="2" data-visibility="2" aria-expanded="false" data-stream-item-id="543542460825" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário para a turma</span></div><div class="Ono85c VvAAB"></div><div jsname="uqYDP" class="QGMq0d Gh0umc kpDQ8 CMmBPd"><div jsaction="JIbuQc:npVELd(IgWJu),sFeBqf(M2UYVd);laiNib:H2nWWd;A56Kbc:BU3G2c;EiG6ec:ZQdNEd; keydown:Hq2uPe" jscontroller="bUQrJd"><div class="QRiHXd"><img aria-hidden="true" alt="" class="a5lbif tkmmwb AI7uec" src="dec2_to_4_files/unnamed_007.jpg" data-atf="false"><div class="a5kY4d cjzpkc-Wvd9Cc QRiHXd yUZA2d"><div class="nxIm7c" jsaction="YqO5N:HRfSZd; keydown:Hq2uPe"><div jsaction="rcuQ6b:rcuQ6b;YFq8g:PqP2y; focus:h06R8" data-role="owner,coteacher,student" data-include-invited="false" jscontroller="r9MpRb" jsname="Ufn6O" jsmodel="LQajt" data-course-id="541227835485"><div class="O98Lj" style=""><div class="bswVrf Lzdwhd-BrZSOd" aria-hidden="true">Adicionar comentário para a turma...</div><div id=":e.t" class="LsqTRb Lzdwhd-AyKMt tgNIJf-Wvd9Cc Yiql6e iTy5c editable" tabindex="0" role="textbox" aria-required="true" aria-multiline="true" aria-label="Adicionar comentário para a turma..." g_editable="true" contenteditable="true"></div></div></div></div><div class="QRiHXd apsLYe "><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db OZ6W0d T8tcPb RDPZE" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="M2UYVd" aria-label="Postar" aria-disabled="true" tabindex="-1" data-tooltip="Postar" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M2 3v18l20-9L2 3zm2 11l9-2-9-2V6.09L17.13 12 4 17.91V14z"></path></svg></span></span></div></div></div></div></div></div></div></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543542307823" class="qhnNic LBlAUc Aopndd TIunU"><div class="n4xnA"><div class="JZicYb QRiHXd"><img class="tnyRnb tkmmwb" aria-hidden="true" src="dec2_to_4_files/unnamed_003.png" data-atf="false"><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Aviso: "a leitura desses textos é necessária…"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Luis Renato Vedovato</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 14 de mar.</span><span aria-hidden="true">14 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543542307823" data-tooltip=" Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 17 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 17 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="false" data-show-bump="true" data-stream-item-id="543542307823" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Oções de aviso"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div><div class="n8F6Jd"><div class="pco8Kc obylVb j70YMc"><span>a leitura desses textos é necessária para o semestre:<br><br>Leitura: <a target="_blank" href="https://revistadedireitodoconsumidor.emnuvens.com.br/rdc/article/view/77">https://revistadedireitodoconsumidor.emnuvens.com.br/rdc/article/view/77</a>&nbsp;<br><br>Leitura: <a target="_blank" href="https://www.portaldeperiodicos.idp.edu.br/direitopublico/article/view/6956">https://www.portaldeperiodicos.idp.edu.br/direitopublico/article/view/6956</a>&nbsp;Felice
 Falivene Baptista , D., Pereira da Silva , L. C. ., &amp; Celeste 
Fonseca , I. (2023). A Natureza Jurídica da Geração Distribuída de 
Energia Elétrica no Brasil. Direito Público, 19(104). <a target="_blank" href="https://doi.org/10.11117/rdp.v19i104.6956">https://doi.org/10.11117/rdp.v19i104.6956</a></span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;wuANJc:.CLIENT;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel="PTCFbe hGbFme BrMJ0e" data-stream-item-id="543542307823" data-is-edit-mode="false" data-filter="0" data-material-parent-id="PTCFbe" data-include-stream-item-materials="true"><div jsname="UYewLd" class="AgzMgb rhFKgc" style="display: none;"><div jsaction="rcuQ6b:rcuQ6b;KtPeHe:rcuQ6b;wuANJc:rcuQ6b" jscontroller="TPuMf" data-parent-id="PTCFbe" jsname="C2Qrw"></div><div class="MlZb9c d3aYgd " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;IKzbTb:Yo3LPb;wuANJc:.CLIENT" jsname="C2Qrw" data-parent-id="PTCFbe" data-mode="7" data-copies-only="false" data-show-originality-analyses="false" data-forms-only="false" data-read-only="false"></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="MlZb9c d3aYgd " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="7" data-material-parent-id="PTCFbe"></div></div></div><div jsname="QkPyvd" class="" style=""></div></div></div></div><div role="region" jsname="EQPzXb" class="s2g3Xd "><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="2" data-visibility="2" aria-expanded="false" data-stream-item-id="543542307823" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário para a turma</span></div><div class="Ono85c VvAAB"></div><div jsname="uqYDP" class="QGMq0d Gh0umc kpDQ8 CMmBPd"><div jsaction="JIbuQc:npVELd(IgWJu),sFeBqf(M2UYVd);laiNib:H2nWWd;A56Kbc:BU3G2c;EiG6ec:ZQdNEd; keydown:Hq2uPe" jscontroller="bUQrJd"><div class="QRiHXd"><img aria-hidden="true" alt="" class="a5lbif tkmmwb AI7uec" src="dec2_to_4_files/unnamed_007.jpg" data-atf="false"><div class="a5kY4d cjzpkc-Wvd9Cc QRiHXd yUZA2d"><div class="nxIm7c" jsaction="YqO5N:HRfSZd; keydown:Hq2uPe"><div jsaction="rcuQ6b:rcuQ6b;YFq8g:PqP2y; focus:h06R8" data-role="owner,coteacher,student" data-include-invited="false" jscontroller="r9MpRb" jsname="Ufn6O" jsmodel="LQajt" data-course-id="541227835485"><div class="O98Lj" style=""><div class="bswVrf Lzdwhd-BrZSOd" aria-hidden="true">Adicionar comentário para a turma...</div><div id=":f.t" class="LsqTRb Lzdwhd-AyKMt tgNIJf-Wvd9Cc Yiql6e iTy5c editable" tabindex="0" role="textbox" aria-required="true" aria-multiline="true" aria-label="Adicionar comentário para a turma..." g_editable="true" contenteditable="true"></div></div></div></div><div class="QRiHXd apsLYe "><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db OZ6W0d T8tcPb RDPZE" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="M2UYVd" aria-label="Postar" aria-disabled="true" tabindex="-1" data-tooltip="Postar" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M2 3v18l20-9L2 3zm2 11l9-2-9-2V6.09L17.13 12 4 17.91V14z"></path></svg></span></span></div></div></div></div></div></div></div></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543539601429" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;Plano da Disciplina&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "Plano da Disciplina"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Luis Renato Vedovato postou um novo material: Plano da Disciplina</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 14 de mar.</span><span aria-hidden="true">14 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543539601429" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 17 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 17 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543539601429" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543539601429"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543539601429"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543511008109" class="qhnNic LBlAUc Aopndd TIunU"><div class="n4xnA"><div class="JZicYb QRiHXd"><img class="tnyRnb tkmmwb" aria-hidden="true" src="dec2_to_4_files/unnamed_004.png" data-atf="false"><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Postada por Giovani Lorenzo Bianchini Dos Santos</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Giovani Lorenzo Bianchini Dos Santos</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 13 de mar.</span><span aria-hidden="true">13 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543511008109" data-tooltip=" Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 16 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 16 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="false" data-show-bump="true" data-stream-item-id="543511008109" class="" id="ow649" __is_owner="true"><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de postagens"><div class="NWlf3e MbhUzd" jsname="ksKsZd" style="top: 26px; left: 13px; width: 40px; height: 40px;"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div><div class="n8F6Jd"><div class="pco8Kc obylVb j70YMc"><span>Eai blz</span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;wuANJc:.CLIENT;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel="PTCFbe hGbFme BrMJ0e" data-stream-item-id="543511008109" data-is-edit-mode="false" data-filter="0" data-material-parent-id="PTCFbe" data-include-stream-item-materials="true"><div jsname="UYewLd" class="AgzMgb rhFKgc" style="display: none;"><div jsaction="rcuQ6b:rcuQ6b;KtPeHe:rcuQ6b;wuANJc:rcuQ6b" jscontroller="TPuMf" data-parent-id="PTCFbe" jsname="C2Qrw"></div><div class="MlZb9c d3aYgd " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;IKzbTb:Yo3LPb;wuANJc:.CLIENT" jsname="C2Qrw" data-parent-id="PTCFbe" data-mode="7" data-copies-only="false" data-show-originality-analyses="false" data-forms-only="false" data-read-only="false"></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="MlZb9c d3aYgd " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="7" data-material-parent-id="PTCFbe"></div></div></div><div jsname="QkPyvd" class="" style=""></div></div></div></div><div role="region" jsname="EQPzXb" class="s2g3Xd "><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="2" data-visibility="2" aria-expanded="false" data-stream-item-id="543511008109" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário para a turma</span></div><div class="Ono85c VvAAB"></div><div jsname="uqYDP" class="QGMq0d Gh0umc kpDQ8 CMmBPd"><div jsaction="JIbuQc:npVELd(IgWJu),sFeBqf(M2UYVd);laiNib:H2nWWd;A56Kbc:BU3G2c;EiG6ec:ZQdNEd; keydown:Hq2uPe" jscontroller="bUQrJd"><div class="QRiHXd"><img aria-hidden="true" alt="" class="a5lbif tkmmwb AI7uec" src="dec2_to_4_files/unnamed_007.jpg" data-atf="false"><div class="a5kY4d cjzpkc-Wvd9Cc QRiHXd yUZA2d"><div class="nxIm7c" jsaction="YqO5N:HRfSZd; keydown:Hq2uPe"><div jsaction="rcuQ6b:rcuQ6b;YFq8g:PqP2y; focus:h06R8" data-role="owner,coteacher,student" data-include-invited="false" jscontroller="r9MpRb" jsname="Ufn6O" jsmodel="LQajt" data-course-id="541227835485"><div class="O98Lj" style=""><div class="bswVrf Lzdwhd-BrZSOd" aria-hidden="true">Adicionar comentário para a turma...</div><div id=":g.t" class="LsqTRb Lzdwhd-AyKMt tgNIJf-Wvd9Cc Yiql6e iTy5c editable" tabindex="0" role="textbox" aria-required="true" aria-multiline="true" aria-label="Adicionar comentário para a turma..." g_editable="true" contenteditable="true"></div></div></div></div><div class="QRiHXd apsLYe "><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db OZ6W0d T8tcPb RDPZE" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="M2UYVd" aria-label="Postar" aria-disabled="true" tabindex="-1" data-tooltip="Postar" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M2 3v18l20-9L2 3zm2 11l9-2-9-2V6.09L17.13 12 4 17.91V14z"></path></svg></span></span></div></div></div></div></div></div></div></div></div><div jsname="ge6pde" class="y9k09d"></div></div></section><div jscontroller="qkFKAf" jsmodel="qjXhl" jsaction="rcuQ6b:ZiN7ye"></div></main></div><div jscontroller="cs6ocd" jsaction="rcuQ6b:npT2md;FttMgb:Qp7hp;qFdNBb:Pb2hxc;Cvbxce:N6n54b;mlnRJb:p5Uonb" style="display: none;" data-wait-for="yidvwe"></div><div jsaction="Cvbxce:ysXIce;qFdNBb:Pb2hxc;uwjiC:xtpvtf;rcuQ6b:npT2md" jscontroller="cpx3"></div><div jsaction="rcuQ6b:OuAj6c;uwjiC:OuAj6c" jscontroller="ZlX84d" id="ow593" __is_owner="true"></div><div jsaction="qFdNBb:Pb2hxc;uwjiC:hDYvKe,bXASFb;FT6KGc:LDHNBf;rcuQ6b:npT2md" jsmodel="xeYtDf" jscontroller="iFgCNe" id="ow570" __is_owner="true"></div></div></div></div><c-data id="c8"></c-data><view-header style="display: none;"><title>Mural</title></view-header></c-wiz><c-wiz c-wiz="" jsrenderer="BZn5fd" class="SSPGKf fXYYpf oCHqfe JwkDRc BIIBbc" jsdata="deferred-c12" data-p="%.@.&quot;NTQxMjM1MjY0NzQ5&quot;]" jscontroller="gQQbc" jsaction="rcuQ6b:rcuQ6b;HO6t5b:PlQWd;gHPzkc:jsAJsc;QmtCl:.CLIENT;qVp5ue:.CLIENT;AE9bOd:.CLIENT;mlnRJb:.CLIENT;uwjiC:.CLIENT" data-node-index="0;0" jsmodel="hc6Ubd PuTOgd;IaLzN;U9kKWe;bYzLLb;lkzLle;" data-ogpc="" data-view-id="ucc-17" data-include-user-lists="true" data-course-states="1" style="visibility: hidden; opacity: 0; position: fixed; inset: -1596px 0px -309px; display: none;" aria-busy="true" data-savescroll="1596" data-savedfocusid="694" aria-hidden="true"><div jsname="a9kxte" class="T4LgNb " style=""><div jsname="qJTHM" class="kFwPee"><div class="xgkURe mhCMAe"></div><div class="xgkURe ECPFEb"></div><div jsaction="rcuQ6b:rcuQ6b" jscontroller="FRimSc"></div><div jsaction="rcuQ6b:rcuQ6b;JIbuQc:hskLsf(ZUkOIc); click:RByGDd(XTYNyb)" role="region" jscontroller="V8Zje" aria-label="Banner informativo" aria-hidden="true"></div><div class="dbEQNc"><div jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:Fmspve(Q7N4Oc);KAD0te:O99HCf" jscontroller="KHqDY" jsmodel="hb3e8b" class="v9TZ3c bFjUmb-Tvm9db"><div class="qyN25"><div class="PFLqgc KFl4Z" style="background-image: url(&quot;https://lh3.googleusercontent.com/hr_crs_themes/AOy-etcoLWshMMuOyuEPi6my1-CGqcB9Xu_JtMHnnqanhyxe6G4JBb0c4t4iCXmTVmGELBHr5m1J3yZjKSy54B4J-1t-DexpdAV-6W6fpizt1pTinEKhdc5iWqk=s1280&quot;);"><div class="VVnuU ra2NV "></div></div><div class="T4tcpe KFl4Z"><h1 class="tNGpbb YrFhrf-ZoZQ1 YVvGBb">G_MC613B_2023S1</h1><div class="qFmcrc z3vRcc-ZoZQ1 YVvGBb"></div></div></div></div><div class="M7zXZd"><aside role="complementary" class="DXLeqd"><div class="CG2qQ dsW6Nd"><div jscontroller="UqV0cb" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b"><div jscontroller="RO1Frf" jsaction="rcuQ6b:rcuQ6b;rKHbQd:r2JIKb;HGIkz:VlevBc;uwjiC:rcuQ6b;JIbuQc:RYcsse(BIFOEb)" class="d4Fe0d LBlAUc NA2Gt" style="display: none;" id="ow724" __is_owner="true"><div class="NGVAIb QRiHXd"><img src="dec2_to_4_files/logo_meet_2020q4_color_1x_web_48dp.png" alt="" aria-hidden="true" class="RponAc" data-atf="false"><span class="asQXV">Meet</span><div class="fPqOAb"></div><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb oxacD" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" aria-label="Opções do link do Meet" aria-disabled="false" tabindex="0" aria-haspopup="true" aria-expanded="false" data-alignright="true"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span><div jsname="xl07Ob" style="display: none;" aria-hidden="true"><div role="menu" tabindex="0" class="JPdR6b hVNH5c" jscontroller="uY3Nvd" jsaction="IpSVtb:TvD9Pc;fEN2Ze:xzS4ub;frq95c:LNeFm;cFpp9e:J9oOtd; click:H8nU8b; mouseup:H8nU8b; keydown:I481le; keypress:Kr2w4b; blur:O22p3e; focus:H8nU8b"><div class="XvhY1d" jsaction="mousedown:p8EH2c; touchstart:p8EH2c"><div class="JAPqpe K0NPx"></div></div></div></div></div></div></div></div><div jscontroller="UqV0cb" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b"></div><div class="d4Fe0d LBlAUc "><div class="WMQb5e" jsmodel="hCpsVc"><h2 class="EZrbnd sxa9Pc">Próximas atividades</h2><div jscontroller="sxyRaf" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;GjA5Zb:rcuQ6b"><div class="lziZub sdDCme"><span class="Y5vSD">Nenhuma atividade para a próxima semana</span><span class="nforOe">Nenhuma atividade para a próxima semana!</span></div><div class="CHJgKd"><div class="VfPpkd-dgl2Hf-ppHlrf-sM5MNb" data-is-touch-wrapper="true"><div class="VfPpkd-LgbsSe VfPpkd-LgbsSe-OWXEXe-dgl2Hf ksBjEc lKxP2d LQeN7 uBUej n42Gr" jscontroller="nKuFpb" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="ksBjEc lKxP2d LQeN7 uBUej n42Gr"><div class="VfPpkd-Jh9lGc"></div><span jsname="V67aGc" class="VfPpkd-vQzf8d" aria-hidden="true">Ver tudo</span><a jsname="hSRGPd" class="WpHeLc VfPpkd-mRLv6 VfPpkd-RLmnJb" href="https://classroom.google.com/a/not-turned-in/NTQxMjM1MjY0NzQ5" aria-label="Ver todas as atividades"></a><div class="VfPpkd-J1Ukfc-LhBDec"></div></div></div></div></div></div></div></div></aside><main class="Sgw65b kdAl3b" jsmodel="uJydvc;I8BbUd;UvJ3Mb;" tabindex="-1" role="main" data-focusid="694"><div jsmodel="NYdJ9b" data-include-stream-item-materials="false" data-stream-item-types="3" data-list-type="5" data-active-filter="1" data-load-all-pages="true"><div jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;oquPK:rcuQ6b;o2F6Cf:if3DMb" jscontroller="s2wDwf"></div></div><section guidedhelpid="streamContentGH" role="section" jsmodel="NYdJ9b" data-include-stream-item-materials="false" data-list-type="3" data-active-filter="2" data-load-all-pages="false"><div jsaction="rcuQ6b:BU4fHd;HO6t5b:BU4fHd;oquPK:E3Ktff;uwjiC:E3Ktff,rcuQ6b;wJx4ze:rcuQ6b;gbLJWc:ZLWxKf;JIbuQc:fyRA7e(idVoDf);gY980b:B9ntFe" jscontroller="yidvwe" id="ow692" __is_owner="true"><div jscontroller="fJcHcd" class="zOtZye LBlAUc GWZ7yf nmFHZb" jsaction="rcuQ6b:rcuQ6b;peFp2d:Fck3Oe;QAK2O:huHkmc;M6YzAd:Bv9PPc"><div class="zTrXGf "><div class="qk0lee QRiHXd VBEdtc-Wvd9Cc" jsaction="click:Fck3Oe" tabindex="0" role="button" guidedhelpid="courseInlineCreatorGH"><div class="U2zcIf"><div jscontroller="tF6Lzd" jsaction="rcuQ6b:rcuQ6b;FZ977b:rcuQ6b"><img class="tkmmwb" jsname="xJzy8c" aria-hidden="true" src="dec2_to_4_files/unnamed_007.jpg" data-atf="false" width="40px" height="40px"></div></div><div class="K6Ovqd">Escreva um aviso para sua turma</div></div><div class="Y5vSD fidHdf" jsaction="JIbuQc:pJN26"><span data-is-tooltip-wrapper="true"><button class="VfPpkd-Bz112c-LgbsSe yHy1rc eT1oJ mN1ivc" jscontroller="soHxf" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc; touchcancel:JMtRjd; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;mlnRJb:fLiPzd" data-idom-class="yHy1rc eT1oJ mN1ivc" jsname="JC5QVe" aria-label="Reutilizar postagem" data-tooltip-enabled="true" data-tooltip-id="tt-c19" guidedhelpid="courseReuseGH"><div jsname="s3Eaab" class="VfPpkd-Bz112c-Jh9lGc"></div><div class="VfPpkd-Bz112c-J1Ukfc-LhBDec"></div><span class="VfPpkd-kBDsod xSP5ic" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M19 5H4v6h2V7h13M5 19h15v-6h-2v4H5"></path><path d="M16.29 10.71l-1.41-1.42L18.17 6l-3.29-3.29 1.41-1.42L21 6zm-8.58 12L3 18l4.71-4.71 1.41 1.42L5.83 18l3.29 3.29z"></path></svg></span></button><div class="EY8ABd-OWXEXe-TAWMXe" role="tooltip" aria-hidden="true" id="tt-c19">Reutilizar postagem</div></span></div></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543535859359" class="qhnNic LBlAUc Aopndd TIunU"><div class="n4xnA"><div class="JZicYb QRiHXd"><img class="tnyRnb tkmmwb" aria-hidden="true" src="dec2_to_4_files/unnamed.png" data-atf="false"><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Aviso: "Horário das monitorias online (via…"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Mateus De Padua Vicente</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 14 de mar.</span><span aria-hidden="true">14 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543535859359" data-tooltip=" Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 17 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta postagem está visível para todos os professores da turma. Ela será permanentemente excluída em 17 dias.</div></div><div><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="false" data-show-bump="true" data-stream-item-id="543535859359" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Oções de aviso"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div><div class="n8F6Jd"><div class="pco8Kc obylVb j70YMc"><span>Horário das monitorias online (via Google Meet):<br><b>Terças-feiras - 15h as 17h</b><br><b>Quintas-feiras - 15h as 17h</b></span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;wuANJc:.CLIENT;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel="PTCFbe hGbFme BrMJ0e" data-stream-item-id="543535859359" data-is-edit-mode="false" data-filter="0" data-material-parent-id="PTCFbe" data-include-stream-item-materials="true"><div jsname="UYewLd" class="AgzMgb rhFKgc" style=""><div jsaction="rcuQ6b:rcuQ6b;KtPeHe:rcuQ6b;wuANJc:rcuQ6b" jscontroller="TPuMf" data-parent-id="PTCFbe" jsname="C2Qrw"></div><div class="MlZb9c d3aYgd " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;IKzbTb:Yo3LPb;wuANJc:.CLIENT" jsname="C2Qrw" data-parent-id="PTCFbe" data-mode="7" data-copies-only="false" data-show-originality-analyses="false" data-forms-only="false" data-read-only="false"><div class="luto0c" data-dom-id="https://meet.google.com/ooo-roex-wdd-0-1-4-https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179-Videochamada com a turma-$$-false-false-false-false-$-$-https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179"><a class="VkhHKd e7EEH nQaZq" target="_blank" aria-label="Anexo: link para https://meet.google.com/ooo-roex-wdd" jsaction="LWntbc" href="https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179" data-focus-id="eTkQDe-https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179" data-attachment-id="https://meet.google.com/ooo-roex-wdd" jsname="HzV7m" data-dom-id="https://meet.google.com/ooo-roex-wdd-0-1-4-https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179-Videochamada com a turma-$$-false-false-false-false-$-$-https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179"><div class="DAnlhb bFjUmb-Wvd9Cc"></div><div class="gM4mlb bFjUmb-Wvd9Cc"></div><div class="rzTfPe xSP5ic "><span class="DPvwYc" aria-hidden="true"></span></div><div class="lIHx8b YVvGBb asQXV ">Videochamada com a turma</div></a><div class="pOf0gc QRiHXd Aopndd M4LFnf" jsname="XgfUnd" data-attachment-id="https://meet.google.com/ooo-roex-wdd" jsaction="JIbuQc:Rsbfue(Rsbfue);"><a class="vwNuXe JkIgWb QRiHXd MymH0d maXJsd" target="_blank" aria-label="Anexo: link para https://meet.google.com/ooo-roex-wdd" jsaction="LWntbc" href="https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179" title="Videochamada com a turma" data-focus-id="hSRGPd-auswjd-https://meet.google.com/ooo-roex-wdd-https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179" data-attachment-id="https://meet.google.com/ooo-roex-wdd"><div class="bxp7vf bHOAdb Niache"><img jsname="q4uQmd" jsaction="error:dyBsCf" class=" " src="dec2_to_4_files/logo_meet_2020q4_color_1x_web_96dp.png" aria-hidden="true" role="presentation" data-mime-type="" data-atf="false"></div><div class="MM30Lb"><div class="A6dC2c QDKOcc VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">Videochamada com a turma</div><div class="cSyPgb WInaFd QRiHXd"><div class="QRiHXd"><div class="kRYv9b YVvGBb">https://meet.google.com/ooo-roex-wdd?authuser=0&amp;hs=179</div></div></div></div></a><div class="ZgfM9 QRiHXd"></div></div></div></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="MlZb9c d3aYgd " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="7" data-material-parent-id="PTCFbe"></div></div></div><div jsname="QkPyvd" class="" style="display: none;"></div></div></div></div><div role="region" jsname="EQPzXb" class="s2g3Xd "><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="2" data-visibility="2" aria-expanded="false" data-stream-item-id="543535859359" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário para a turma</span></div><div class="Ono85c VvAAB"></div><div jsname="uqYDP" class="QGMq0d Gh0umc kpDQ8 CMmBPd"><div jsaction="JIbuQc:npVELd(IgWJu),sFeBqf(M2UYVd);laiNib:H2nWWd;A56Kbc:BU3G2c;EiG6ec:ZQdNEd; keydown:Hq2uPe" jscontroller="bUQrJd"><div class="QRiHXd"><img aria-hidden="true" alt="" class="a5lbif tkmmwb AI7uec" src="dec2_to_4_files/unnamed_007.jpg" data-atf="false"><div class="a5kY4d cjzpkc-Wvd9Cc QRiHXd yUZA2d"><div class="nxIm7c" jsaction="YqO5N:HRfSZd; keydown:Hq2uPe"><div jsaction="rcuQ6b:rcuQ6b;YFq8g:PqP2y; focus:h06R8" data-role="owner,coteacher,student" data-include-invited="false" jscontroller="r9MpRb" jsname="Ufn6O" jsmodel="LQajt" data-course-id="541235264749"><div class="O98Lj" style=""><div class="bswVrf Lzdwhd-BrZSOd" aria-hidden="true">Adicionar comentário para a turma...</div><div id=":h.t" class="LsqTRb Lzdwhd-AyKMt tgNIJf-Wvd9Cc Yiql6e iTy5c editable" tabindex="0" role="textbox" aria-required="true" aria-multiline="true" aria-label="Adicionar comentário para a turma..." g_editable="true" contenteditable="true"></div></div></div></div><div class="QRiHXd apsLYe "><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db OZ6W0d T8tcPb RDPZE" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="M2UYVd" aria-label="Postar" aria-disabled="true" tabindex="-1" data-tooltip="Postar" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M2 3v18l20-9L2 3zm2 11l9-2-9-2V6.09L17.13 12 4 17.91V14z"></path></svg></span></span></div></div></div></div></div></div></div></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543338621102" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;DATAS DE ENTREGA DOS LABORATÓRIOS&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "DATAS DE ENTREGA DOS LABORATÓRIOS"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou um novo material: DATAS DE ENTREGA DOS LABORATÓRIOS</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543338621102" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 11 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 11 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543338621102" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543338621102"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543338621102"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543338359528" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;MC602 - TEORIA CIRCUITOS LÓGICOS&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "MC602 - TEORIA CIRCUITOS LÓGICOS"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou um novo material: MC602 - TEORIA CIRCUITOS LÓGICOS</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543338359528" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 11 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 11 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543338359528" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543338359528"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543338359528"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303561243" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB12&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB12"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB12</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303561243" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303561243" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303561243"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303561243"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303471225" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB11&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB11"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB11</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303471225" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303471225" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303471225"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303471225"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303370649" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB10&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB10"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB10</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303370649" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303370649" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303370649"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303370649"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303497207" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB09&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB09"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB09</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303497207" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303497207" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303497207"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303497207"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303493100" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB08&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB08"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB08</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303493100" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303493100" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303493100"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303493100"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303423666" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB07&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB07"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB07</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303423666" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303423666" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303423666"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303423666"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303465543" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB06&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB06"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB06</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303465543" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303465543" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303465543"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303465543"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303377608" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB05&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB05"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB05</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303377608" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303377608" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303377608"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543303377608"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="563082264962" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB04&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB04"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB04</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-563082264962" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="563082264962" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="563082264962"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|563082264962"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303401379" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB03&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB03"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB03</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303401379" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303401379" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303401379"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="false" data-focus-id="LPEWg|543303401379"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"><span class="VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">2 comentários da turma</span></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303423454" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB02&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB02"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB02</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303423454" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 11 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 11 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303423454" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303423454"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="false" data-focus-id="LPEWg|543303423454"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"><span class="VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">2 comentários da turma</span></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543303407617" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Atividade: &quot;LAB01&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Atividade: "LAB01"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou uma nova atividade: LAB01</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 8 de mar.</span><span aria-hidden="true">8 de mar.</span>&nbsp;Editado às 21 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543303407617" data-tooltip=" Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Esta atividade está visível para todos os professores da turma. Ela será permanentemente excluída em 24 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543303407617" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543303407617"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="false" data-focus-id="LPEWg|543303407617"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"><span class="VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc"> 1 comentário para a turma</span></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543129813778" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;DE1 SoC BOARD&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "DE1 SoC BOARD"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou um novo material: DE1 SoC BOARD</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 3 de mar.</span><span aria-hidden="true">3 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543129813778" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543129813778" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543129813778"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543129813778"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543130420311" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;SLIDES DE AULAS&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "SLIDES DE AULAS"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou um novo material: SLIDES DE AULAS</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 3 de mar.</span><span aria-hidden="true">3 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543130420311" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543130420311" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543130420311"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543130420311"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543129452865" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;DATA DE ENTREGA DOS LABORATÓRIOS&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "DATA DE ENTREGA DOS LABORATÓRIOS"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou um novo material: DATA DE ENTREGA DOS LABORATÓRIOS</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 3 de mar.</span><span aria-hidden="true">3 de mar.</span>&nbsp;Editado às 8 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543129452865" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 11 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 11 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543129452865" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543129452865"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543129452865"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543129518247" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;PROGRAMA DISCIPLINA MC613 TURMA B&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "PROGRAMA DISCIPLINA MC613 TURMA B"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou um novo material: PROGRAMA DISCIPLINA MC613 TURMA B</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 3 de mar.</span><span aria-hidden="true">3 de mar.</span><span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543129518247" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543129518247" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543129518247"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543129518247"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsmodel="PTCFbe" data-include-stream-item-materials="false" data-stream-item-id="543128966291" jsaction="click:YdzvGf" class="qhnNic LBlAUc Aopndd TIunU ZoT1D idtp4e DkDwHe"><div class="n4xnA"><div class="JZicYb QRiHXd"><div class="PazDv" jsname="rQC7Ie" tabindex="0" role="link" aria-label="Material: &quot;AULAS GRAVADAS -  LINKS&quot;"></div><div class="bxp7vf bFjUmb-Wvd9Cc m1PbN qJJSvb vUBwW"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M18 2H6c-1.1 0-2 .9-2 2v16c0 1.1.9 2 2 2h12c1.1 0 2-.9 2-2V4c0-1.1-.9-2-2-2zm0 18H6V4h2v8l2.5-1.5L13 12V4h5v16z"></path></svg></div><div class="GQW44b"><div class="lziZub tLDEHd"><h2><span class="PazDv">Material: "AULAS GRAVADAS -  LINKS"</span></h2><div class="QRiHXd"><span class="YVvGBb asQXV">Ricardo Pannain postou um novo material: AULAS GRAVADAS -  LINKS</span></div></div><span class="IMvYId dDKhVc YVvGBb"><span class="PazDv">Criado em: 3 de mar.</span><span aria-hidden="true">3 de mar.</span>&nbsp;Editado às 3 de mar.<span class="IMvYId P354se"> – Excluído</span></span></div><div class="Nmpzvc"></div><div jscontroller="By0w6" jsaction="mouseover:eGiyHb; click:eGiyHb; focus:eGiyHb; touchstart:eGiyHb" role="tooltip" tabindex="0" data-focus-id="IlqLNc-543128966291" data-tooltip=" Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias." class="a7OWub  JEf8lc P354se"><span class="xSP5ic "><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M11 18h2v-2h-2v2zm1-16C6.48 2 2 6.48 2 12s4.48 10 10 10 10-4.48 10-10S17.52 2 12 2zm0 18c-4.41 0-8-3.59-8-8s3.59-8 8-8 8 3.59 8 8-3.59 8-8 8zm0-14c-2.21 0-4 1.79-4 4h2c0-1.1.9-2 2-2s2 .9 2 2c0 2-3 1.75-3 5h2c0-2.25 3-2.5 3-5 0-2.21-1.79-4-4-4z"></path></svg></span><div class="PazDv" jsname="bOjMyf"> Este material está visível para todos os professores desta turma. Ele será excluído permanentemente em 6 dias.</div></div><div data-guided-help-id="streamItemActionMenuGH"><div class="kpDQ8 qZsscc"><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;oquPK:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:N6Gb7c" data-hide-copy-link="false" data-hide-delete="true" data-show-bump="true" data-stream-item-id="543128966291" class=""><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções do material"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div></div></div></div><div class="BoJUHd" jsmodel="xvu37b" jsaction="rg93rb" data-type="2" data-visibility="2" data-stream-item-id="543128966291"><a class="onkcGd JX1kZ VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc" target="_self" jsname="HeH4ab" aria-hidden="true" data-focus-id="LPEWg|543128966291"><div jscontroller="QdwYy" jsaction="rcuQ6b:.rcuQ6b;Ts0WYd:.rcuQ6b" data-comment-type="2" data-hide-if-zero="true" data-ancestor-selector=".JX1kZ" class="QSmq3c ZNE4y"></div></a></div></div><div jsname="ge6pde" class="y9k09d"></div></div></section><div jscontroller="qkFKAf" jsmodel="qjXhl" jsaction="rcuQ6b:ZiN7ye"></div></main></div><div jscontroller="cs6ocd" jsaction="rcuQ6b:npT2md;FttMgb:Qp7hp;qFdNBb:Pb2hxc;Cvbxce:N6n54b;mlnRJb:p5Uonb" style="display: none;" data-wait-for="yidvwe"></div><div jsaction="Cvbxce:ysXIce;qFdNBb:Pb2hxc;uwjiC:xtpvtf;rcuQ6b:npT2md" jscontroller="cpx3"></div><div jsaction="rcuQ6b:OuAj6c;uwjiC:OuAj6c" jscontroller="ZlX84d" id="ow714" __is_owner="true"></div><div jsaction="qFdNBb:Pb2hxc;uwjiC:hDYvKe,bXASFb;FT6KGc:LDHNBf;rcuQ6b:npT2md" jsmodel="xeYtDf" jscontroller="iFgCNe" id="ow691" __is_owner="true"></div></div></div></div><c-data id="c12"></c-data><view-header style="display: none;"><title>Mural</title></view-header></c-wiz><c-wiz c-wiz="" jsrenderer="eTaVhe" class="SSPGKf fXYYpf JwkDRc oCHqfe BIIBbc" jsdata="deferred-c18" data-p="%.@.&quot;NTQxMjM1MjY0NzQ5&quot;,&quot;a&quot;,&quot;NTQzMzAzNDA3NjE3&quot;]" jscontroller="gQQbc" jsaction="rcuQ6b:rcuQ6b;HO6t5b:PlQWd;gHPzkc:jsAJsc;QmtCl:.CLIENT;qVp5ue:.CLIENT;AE9bOd:.CLIENT;mlnRJb:.CLIENT;uwjiC:.CLIENT;wuANJc:.CLIENT;voP7ud:.CLIENT" data-node-index="0;0" jsmodel="hc6Ubd PuTOgd;IaLzN;U9kKWe;bYzLLb;PTCFbe;dSSknb;lkzLle;r5HSpf;" data-ogpc="" data-view-id="ucc-18" data-include-user-lists="true" data-include-stream-item-materials="false" data-without-stream-item-materials="" data-submission-id="2" data-force-create="true" data-include-submission-materials="true" style="visibility: hidden; opacity: 0; position: fixed; inset: 0px 0px 137.5px; display: none;" aria-busy="true" data-savescroll="0" data-savedfocusid="984" aria-hidden="true"><div jsname="a9kxte" class="T4LgNb "><div jsname="qJTHM" class="kFwPee"><div class="xgkURe mhCMAe"></div><div class="xgkURe ECPFEb"></div><div jsaction="rcuQ6b:rcuQ6b" jscontroller="FRimSc"></div><div jscontroller="UqV0cb" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b"><div jscontroller="cs6ocd" jsaction="rcuQ6b:npT2md;FttMgb:Qp7hp;qFdNBb:Pb2hxc;Cvbxce:N6n54b;mlnRJb:p5Uonb" style="display: none;" data-wait-for="QlRoyd"></div><div class="fJ1Vac"><div class="P47N4e vUBwW m1PbN bFjUmb-Wvd9Cc pOf0gc"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="EE538" role="main"><div jscontroller="QlRoyd" jsmodel="I8BbUd;UvJ3Mb;uJydvc;xeYtDf;" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;wJx4ze:rcuQ6b"><div class="nl5VRd ypv4re"><div class="N5dSp"><h1 class="fOvfyc B7SYid VnOHwf-Tvm9db"><span style="white-space: pre-wrap;">LAB01</span></h1><div class="Nmpzvc"></div><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:yG0upc" data-hide-copy-link="false" data-hide-delete="false" data-stream-item-id="543303407617" class="I0naMd"><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb wwnMtb oxacD" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div><div class="rec5Nb cSyPgb QRiHXd"><div class="YVvGBb">Ricardo Pannain</div><div class="DwLQSc" aria-hidden="true">•</div><div class="YVvGBb">8 de mar.&nbsp;Editado às 21 de mar.</div></div><div class="W4hhKd"><div class="CzuI5c asQXV QRiHXd"><div class="YVvGBb"><div jsaction="rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b" jscontroller="teDhve"><div aria-hidden="true">0,28<span class="AgnJoc">/1</span></div><div class="PazDv">0,28 ponto de 1 possíveis</div></div></div></div><div class="asQXV hnID5d"></div></div><div class="Wa3mee nQaZq"><div jscontroller="IGT0cf" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;JIbuQc:Yh7j1c(PlbUX)" jsmodel="xvu37b" data-type="2" data-visibility="2" guidedhelpid="commentsdialogGH" class=" LhPqk" data-with-icon="true" data-show-add-comments-link="true"><div role="button" class="uArJ5e cd29Sd UQuaGc kCyAyd oxacD" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;" jsshadow="" jsname="PlbUX" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue cd29Sd"><span class="E6FpNe Ce1Y1c"><svg width="24" height="24" viewBox="0 0 24 24" focusable="false" class=" NMm5M hhikbc"><path d="M21.99 4c0-1.1-.89-2-1.99-2H4c-1.1 0-2 .9-2 2v12c0 1.1.9 2 2 2h14l4 4-.01-18zM4 16V4h16v12H4z"></path><path d="M6 12h12v2H6zm0-3h12v2H6zm0-3h12v2H6z"></path></svg></span><span class="NPEfkd RveJvd snByac"> 1 comentário para a turma</span></span></div></div></div></div></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;wuANJc:.CLIENT;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel="PTCFbe hGbFme BrMJ0e" data-is-edit-mode="false" data-filter="0" data-material-parent-id="PTCFbe" data-include-stream-item-materials="true"><div jsname="UYewLd" class="AgzMgb hjqfGd" style=""><div class="MlZb9c xLFtvb " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;IKzbTb:Yo3LPb;wuANJc:.CLIENT" jsname="C2Qrw" data-parent-id="PTCFbe" data-mode="1" data-copies-only="false" data-show-originality-analyses="false" data-forms-only="false" data-read-only="false"><div data-dom-id="1-Yrut9yc__AHCb0tRLe6Ct9jV0NioUXU-0-1-2-PDF-lab01_v2023.1.pdf-$2-false-false-false-false-$-$-https://drive.google.com/file/d/1-Yrut9yc__AHCb0tRLe6Ct9jV0NioUXU/view?usp=drive_web&amp;authuser=0" class="t2wIBc"><div class="r0VQac QRiHXd Aopndd " jsname="HzV7m" jsaction="JIbuQc:Rsbfue(Rsbfue);"><a class="vwNuXe JkIgWb QRiHXd MymH0d maXJsd" target="_blank" aria-label="Anexo: PDF: lab01_v2023.1.pdf" jsaction="LWntbc" href="https://drive.google.com/file/d/1-Yrut9yc__AHCb0tRLe6Ct9jV0NioUXU/view?usp=drive_web&amp;authuser=0" title="lab01_v2023.1.pdf" data-focus-id="hSRGPd-auswjd-1-Yrut9yc__AHCb0tRLe6Ct9jV0NioUXU-https://drive.google.com/file/d/1-Yrut9yc__AHCb0tRLe6Ct9jV0NioUXU/view?usp=drive_web&amp;authuser=0" data-attachment-id="1-Yrut9yc__AHCb0tRLe6Ct9jV0NioUXU" data-focusid="984"><div class="bxp7vf bHOAdb Niache"><img jsname="q4uQmd" jsaction="error:dyBsCf" class=" " src="dec2_to_4_files/lab01_v2023.1.pdf.png" aria-hidden="true" role="presentation" data-mime-type="application/pdf" data-atf="false"></div><div class="MM30Lb"><div class="A6dC2c QDKOcc VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">lab01_v2023.1.pdf</div><div class="cSyPgb WInaFd QRiHXd"><div class="QRiHXd"><div class="kRYv9b YVvGBb">PDF</div></div></div></div></a><div class="ZgfM9 QRiHXd"></div></div></div></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="MlZb9c xLFtvb " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="1" data-material-parent-id="PTCFbe"></div></div></div><div jsname="QkPyvd" class="" style="display: none;"></div></div><div jsmodel="WuwnAd;jmgIWd;" jscontroller="F37rhb" jsaction="rcuQ6b:rcuQ6b;LSbPUe:rcuQ6b;voP7ud:rcuQ6b" data-course-id="541235264749" class="Z3wmOd lLBkgb" data-allow-rubric-scoring="false"></div><div class="smtc7c"><div class="GWZ7yf AJFihd LBlAUc YkTkoe"><div class="Dy8Cxc QRiHXd"><span class="z3vRcc">Seus trabalhos<div jscontroller="FQo2Xb" jsaction="rcuQ6b:hDYvKe;voP7ud:hDYvKe;qFdNBb:Pb2hxc"></div></span><span class="asQXV"><span jsaction="rcuQ6b:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;uwjiC:rcuQ6b" jscontroller="o5ZA8b" class="UhYXkc KI1A1e ZnNi8e" data-submission-id="2" data-render-simple-labels="true"><span class="u7S8tc YVvGBb">Com nota</span><span class="E70Hue neggzd" aria-hidden="true">Estigfend</span></span></span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel=" hGbFme BrMJ0e" data-is-edit-mode="false" data-filter="1" data-material-parent-id="2"><div jsname="UYewLd" class="AgzMgb " style="display: none;"><div jscontroller="KqB22e" jsmodel="I8BbUd;PTCFbe;" data-include-stream-item-materials="true" jsaction="rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;mbUMkc:rcuQ6b;IKzbTb:Yo3LPb;wJx4ze:rcuQ6b" jsname="C2Qrw" class="CG2qQ P2wHlc" style="display: none;"></div><div class="JY4wBc MlZb9c " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;IKzbTb:Yo3LPb" jsname="C2Qrw" data-parent-id="2" data-mode="6" data-copies-only="false" data-show-originality-analyses="true" data-forms-only="false" data-read-only="false"></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="JY4wBc MlZb9c " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="6" data-material-parent-id="2"></div></div></div><div jsname="QkPyvd" class="Jp15We tLDEHd B2pRjc" style="">Nenhum trabalho anexado</div><div class="IPGLSb"><div class="QRiHXd J2Cevf" guidedhelpid="submissionManager"><div jsaction="rcuQ6b:rcuQ6b;ln5gI:rcuQ6b;RwVyRc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:rcuQ6b;LEpEAf:qRU3cb" jscontroller="PykWJd" jsmodel="AKq4rd" data-user-id="30751363934" data-attach-actions-control-type="3" data-parent-id="2" class="TDK0Zb CG2qQ cYYbdd"><div jsshadow="" role="button" class="U26fgb REtOWc cd29Sd p0oLxb BEAGS" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" aria-disabled="false" tabindex="0" aria-haspopup="true" aria-expanded="false" guidedhelpid="addOrCreateMaterial" data-menu-type="3" id="ow916" __is_owner="true"><div class="bnqxkd MbhUzd" jsname="ksKsZd"></div><div class="GJYBjd CeoRYc" aria-hidden="true"></div><span jsslot="" class="GcVcmc Fxmcue cd29Sd"><span class="lRRqZc Ce1Y1c"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="a7AG0 NMm5M"><path d="M20 13h-7v7h-2v-7H4v-2h7V4h2v7h7v2z"></path></svg></span><span class="RdyDwe snByac">Adicionar ou criar</span></span></div></div></div><div jscontroller="Glz2Ld" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;JIbuQc:f2nbFb" data-submission-id="2"></div><div jscontroller="krEUN" jsaction="JIbuQc:sFeBqf(sFeBqf),ReqGfd(ReqGfd);rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;nK3Vsc:rcuQ6b;ZQcBrc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:Yo3LPb;R6l5Vd:UApqrc;LNlWBf:IyXkod" class="CG2qQ kg6ice"><div jsshadow="" role="button" class="uArJ5e TuHiFd UQuaGc Y5sE8d" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="sFeBqf" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Enviar novamente</span></span></div></div></div></div><div jscontroller="cTy1kf" jsmodel="I8BbUd" jsaction="rcuQ6b:TZH2db;wuANJc:TZH2db;voP7ud:TZH2db;wJx4ze:TZH2db"></div></div><div class="GWZ7yf m8BrFf LBlAUc YkTkoe" guidedhelpid="submissionPrivateComments"><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="3" data-visibility="1" data-submission-id="30751363934" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;wuANJc:lswmYb;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário particular</span></div><div class="amzDAb"><div class="QxGMXc asQXV QRiHXd"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Comentários particulares</span></div><div jsshadow="" role="button" class="uArJ5e UQuaGc kCyAyd l3F1ye Epqnjf xAiME" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="zPiFrf" aria-label="Adicionar comentário para Ricardo Pannain" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Adicionar comentário para Ricardo Pannain</span></span></div></div><div class="Ono85c VvAAB"></div></div></div></div><div class="pOf0gc"><div class="eqqrO"><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="2" data-visibility="2" class="PeGHgb Q8U8uc" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="VYv8If QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">1 comentário para a turma</span></div><div class="amzDAb"><div class="lq45g asQXV QRiHXd"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">Comentários da turma</span></div></div><div class="ruTJle VvAAB"><div class="dZVZab"><div jsaction="ym8qYd:u4pxTb" jscontroller="dvgIje" class="wJ76ge TIunU"><div class="QRiHXd pMq3Db"><img class="WqfsMd tkmmwb" aria-hidden="true" alt="" src="dec2_to_4_files/unnamed_003.jpg" data-atf="false"><div class="G0rp"><div class="YU7iib"><div><a class="gJItbc asQXV" aria-label="Comentário postado por Ricardo Pannain">Ricardo Pannain</a><span class="T8rTjd">21 de mar.</span></div><div class="thiSD Gh0umc" jsaction="JIbuQc:pODwA(IgWJu)"><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db L8jEMd CMmBPd oxacD qk5dFc kpDQ8" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="IgWJu" aria-label="Responder" tabindex="0" data-tooltip="Responder a este comentário" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M16 10H6.83L9 7.83l1.41-1.41L9 5l-6 6 6 6 1.41-1.41L9 14.17 6.83 12H16c1.65 0 3 1.35 3 3v4h2v-4c0-2.76-2.24-5-5-5z"></path></svg></span></span></div><div class="KYmC8d kpDQ8 CG2qQ"><div jscontroller="RrRSXd" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b" jsmodel="I8BbUd" data-comment-id="543779294004"></div></div></div></div><div class="VSWCL tLDEHd"><span style="white-space: pre-wrap;">NOTA MÁXIMA DO LAB01 É 0,28</span></div></div></div></div></div></div><div jsname="uqYDP" class="XNP4U Gh0umc kpDQ8 CMmBPd"><div jsaction="JIbuQc:npVELd(IgWJu),sFeBqf(M2UYVd);laiNib:H2nWWd;A56Kbc:BU3G2c;EiG6ec:ZQdNEd; keydown:Hq2uPe" jscontroller="bUQrJd"><div class="QRiHXd"><img aria-hidden="true" alt="" class="a5lbif tkmmwb AI7uec" src="dec2_to_4_files/unnamed_007.jpg" data-atf="false"><div class="a5kY4d cjzpkc-Wvd9Cc QRiHXd yUZA2d"><div class="nxIm7c" jsaction="YqO5N:HRfSZd; keydown:Hq2uPe"><div jsaction="rcuQ6b:rcuQ6b;YFq8g:PqP2y; focus:h06R8" data-role="owner,coteacher,student" data-include-invited="false" jscontroller="r9MpRb" jsname="Ufn6O" jsmodel="LQajt" data-course-id="541235264749"><div class="O98Lj" style=""><div class="bswVrf Lzdwhd-BrZSOd" aria-hidden="true">Adicionar comentário para a turma...</div><div id=":i.t" class="LsqTRb Lzdwhd-AyKMt tgNIJf-Wvd9Cc Yiql6e iTy5c editable" tabindex="0" role="textbox" aria-required="true" aria-multiline="true" aria-label="Adicionar comentário para a turma..." g_editable="true" contenteditable="true"></div></div></div></div><div class="QRiHXd apsLYe "><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db OZ6W0d T8tcPb RDPZE" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="M2UYVd" aria-label="Postar" aria-disabled="true" tabindex="-1" data-tooltip="Postar" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M2 3v18l20-9L2 3zm2 11l9-2-9-2V6.09L17.13 12 4 17.91V14z"></path></svg></span></span></div></div></div></div></div></div></div></div></div></div><aside class="asCVDb BiaLW" role="complementary"><div class="GWZ7yf AJFihd LBlAUc YkTkoe"><div class="Dy8Cxc QRiHXd"><span class="z3vRcc">Seus trabalhos<div jscontroller="FQo2Xb" jsaction="rcuQ6b:hDYvKe;voP7ud:hDYvKe;qFdNBb:Pb2hxc"></div></span><span class="asQXV"><span jsaction="rcuQ6b:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;uwjiC:rcuQ6b" jscontroller="o5ZA8b" class="UhYXkc KI1A1e ZnNi8e" data-submission-id="2" data-render-simple-labels="true"><span class="u7S8tc YVvGBb">Com nota</span><span class="E70Hue neggzd" aria-hidden="true">Estigfend</span></span></span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel=" hGbFme BrMJ0e" data-is-edit-mode="false" data-filter="1" data-material-parent-id="2"><div jsname="UYewLd" class="AgzMgb " style="display: none;"><div jscontroller="KqB22e" jsmodel="I8BbUd;PTCFbe;" data-include-stream-item-materials="true" jsaction="rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;mbUMkc:rcuQ6b;IKzbTb:Yo3LPb;wJx4ze:rcuQ6b" jsname="C2Qrw" class="CG2qQ P2wHlc" style="display: none;"></div><div class="JY4wBc MlZb9c " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;IKzbTb:Yo3LPb" jsname="C2Qrw" data-parent-id="2" data-mode="6" data-copies-only="false" data-show-originality-analyses="true" data-forms-only="false" data-read-only="false"></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="JY4wBc MlZb9c " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="6" data-material-parent-id="2"></div></div></div><div jsname="QkPyvd" class="Jp15We tLDEHd B2pRjc" style="">Nenhum trabalho anexado</div><div class="IPGLSb"><div class="QRiHXd J2Cevf" guidedhelpid="submissionManager"><div jsaction="rcuQ6b:rcuQ6b;ln5gI:rcuQ6b;RwVyRc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:rcuQ6b;LEpEAf:qRU3cb" jscontroller="PykWJd" jsmodel="AKq4rd" data-user-id="30751363934" data-attach-actions-control-type="3" data-parent-id="2" class="TDK0Zb CG2qQ cYYbdd"><div jsshadow="" role="button" class="U26fgb REtOWc cd29Sd p0oLxb BEAGS" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" aria-disabled="false" tabindex="0" aria-haspopup="true" aria-expanded="false" guidedhelpid="addOrCreateMaterial" data-menu-type="3"><div class="bnqxkd MbhUzd" jsname="ksKsZd"></div><div class="GJYBjd CeoRYc" aria-hidden="true"></div><span jsslot="" class="GcVcmc Fxmcue cd29Sd"><span class="lRRqZc Ce1Y1c"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="a7AG0 NMm5M"><path d="M20 13h-7v7h-2v-7H4v-2h7V4h2v7h7v2z"></path></svg></span><span class="RdyDwe snByac">Adicionar ou criar</span></span><div jsname="xl07Ob" style="display: none;" aria-hidden="true"><div role="menu" tabindex="0" class="JPdR6b e5Emjc hVNH5c" jscontroller="uY3Nvd" jsaction="IpSVtb:TvD9Pc;fEN2Ze:xzS4ub;frq95c:LNeFm;cFpp9e:J9oOtd; click:H8nU8b; mouseup:H8nU8b; keydown:I481le; keypress:Kr2w4b; blur:O22p3e; focus:H8nU8b"><div class="XvhY1d" jsaction="mousedown:p8EH2c; touchstart:p8EH2c"><div class="JAPqpe K0NPx"><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Google Drive" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg enable-background="new 0 0 24 24" focusable="false" height="24" viewBox="0 0 24 24" width="24" class="zAg7wc xSP5ic NMm5M"><rect fill="none" height="24" width="24"></rect><path d="M14.35,2.5h-4.7c-0.71,0-1.37,0.38-1.73,0.99L1.58,14.4c-0.36,0.62-0.36,1.38-0.01,2l2.35,4.09c0.36,0.62,1.02,1,1.73,1 h12.68c0.72,0,1.38-0.38,1.73-1l2.35-4.09c0.36-0.62,0.35-1.38-0.01-2L16.08,3.49C15.72,2.88,15.06,2.5,14.35,2.5z M18.34,19.5H5.66 l-2.35-4.09L9.65,4.5h4.7l6.34,10.91L18.34,19.5z M12.9,7.75h-1.8l-4.58,7.98L7.25,17h9.5l0.73-1.27L12.9,7.75z M9.25,15L12,10.2 l2.75,4.8H9.25z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:pau0Hb" data-type="2"><div class="jO7h3c">Google Drive</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Link" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="zAg7wc xSP5ic NMm5M"><path d="M3.9 12c0-1.71 1.39-3.1 3.1-3.1h4V7H7c-2.76 0-5 2.24-5 5s2.24 5 5 5h4v-1.9H7c-1.71 0-3.1-1.39-3.1-3.1zM8 13h8v-2H8v2zm9-6h-4v1.9h4c1.71 0 3.1 1.39 3.1 3.1s-1.39 3.1-3.1 3.1h-4V17h4c2.76 0 5-2.24 5-5s-2.24-5-5-5z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:VORrnc"><div class="jO7h3c">Link</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Arquivo" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="zAg7wc xSP5ic NMm5M"><path d="M15.5 6v10.5c0 2.21-1.79 4-4 4s-4-1.79-4-4V6a2.5 2.5 0 0 1 5 0v9.5c0 .55-.45 1-1 1s-1-.45-1-1V6H9v9.5a2.5 2.5 0 0 0 5 0V6c0-2.21-1.79-4-4-4S6 3.79 6 6v10.5c0 3.04 2.46 5.5 5.5 5.5s5.5-2.46 5.5-5.5V6h-1.5z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:pau0Hb" data-type="1"><div class="jO7h3c">Arquivo</div></div></span><div role="separator" aria-hidden="true" class="kCtYwe"></div><h3 class="mMfeif ubvFYc dDKhVc-Wvd9Cc">Criar novo</h3><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Documentos" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="XxyAsb"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="1"><div class="jO7h3c">Documentos</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Apresentações" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="qurv4d"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="3"><div class="jO7h3c">Apresentações</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Planilhas" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="teCq2b"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="2"><div class="jO7h3c">Planilhas</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Desenhos" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="O1YELb"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="6"><div class="jO7h3c">Desenhos</div></div></span></div></div></div></div></div></div></div><div jscontroller="Glz2Ld" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;JIbuQc:f2nbFb" data-submission-id="2"></div><div jscontroller="krEUN" jsaction="JIbuQc:sFeBqf(sFeBqf),ReqGfd(ReqGfd);rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;nK3Vsc:rcuQ6b;ZQcBrc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:Yo3LPb;R6l5Vd:UApqrc;LNlWBf:IyXkod" class="CG2qQ kg6ice"><div jsshadow="" role="button" class="uArJ5e TuHiFd UQuaGc Y5sE8d" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="sFeBqf" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Enviar novamente</span></span></div></div></div></div><div jscontroller="cTy1kf" jsmodel="I8BbUd" jsaction="rcuQ6b:TZH2db;wuANJc:TZH2db;voP7ud:TZH2db;wJx4ze:TZH2db"></div></div><div class="GWZ7yf m8BrFf LBlAUc YkTkoe" guidedhelpid="submissionPrivateComments"><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="3" data-visibility="1" data-submission-id="30751363934" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;wuANJc:lswmYb;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário particular</span></div><div class="amzDAb"><div class="QxGMXc asQXV QRiHXd"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Comentários particulares</span></div><div jsshadow="" role="button" class="uArJ5e UQuaGc kCyAyd l3F1ye Epqnjf xAiME" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="zPiFrf" aria-label="Adicionar comentário para Ricardo Pannain" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Adicionar comentário para Ricardo Pannain</span></span></div></div><div class="Ono85c VvAAB"></div></div></div></aside></div></div><div jscontroller="rFwfKe" jsaction="qFdNBb:Pb2hxc;pN3Oaf:n3lXYe;uwjiC:T0iadd;wuANJc:T0iadd;voP7ud:T0iadd"></div><div jscontroller="BbOAsf" jsmodel="PTCFbe;" jsaction="qFdNBb:Pb2hxc;Cvbxce:ysXIce;pN3Oaf:n3lXYe;wuANJc:hDYvKe,T0iadd;ywGDo:hDYvKe;rcuQ6b:npT2md" data-include-stream-item-materials="true" data-with-stream-item-materials=""></div><div jsaction="Cvbxce:ysXIce;qFdNBb:Pb2hxc;uwjiC:xtpvtf;rcuQ6b:npT2md" jscontroller="cpx3"></div><div jsaction="rcuQ6b:OuAj6c;uwjiC:OuAj6c" jscontroller="ZlX84d" id="ow893" __is_owner="true"></div></div></div><c-data id="c18"></c-data><view-header style="display: none;"><title>Detalhes da atividade</title></view-header></c-wiz><div jscontroller="HmEm0" jsaction="BfpAHf:TCTP9d;Nwyqre:DsZxZc; transitionend:e204de;O0KOhf:.CLIENT;SemCgb:.CLIENT" id="tt-i1-visible-label" class="VfPpkd-suEOdc EY8ABd" aria-hidden="true"><div class="VfPpkd-z59Tgd VfPpkd-z59Tgd-OiiCO"><span class="VfPpkd-A3KfFd">Menu principal</span></div></div><c-wiz c-wiz="" jsrenderer="eTaVhe" class="SSPGKf fXYYpf" jsdata="deferred-c20" data-p="%.@.&quot;NTQxMjM1MjY0NzQ5&quot;,&quot;a&quot;,&quot;NTQzMzAzNDAxMzc5&quot;]" jscontroller="gQQbc" jsaction="rcuQ6b:rcuQ6b;HO6t5b:PlQWd;gHPzkc:jsAJsc;QmtCl:.CLIENT;qVp5ue:.CLIENT;AE9bOd:.CLIENT;mlnRJb:.CLIENT;uwjiC:.CLIENT;wuANJc:.CLIENT;voP7ud:.CLIENT" data-node-index="0;0" jsmodel="hc6Ubd PuTOgd;IaLzN;U9kKWe;bYzLLb;PTCFbe;dSSknb;lkzLle;r5HSpf;" data-ogpc="" data-view-id="ucc-19" data-include-user-lists="true" data-include-stream-item-materials="false" data-without-stream-item-materials="" data-submission-id="2" data-force-create="true" data-include-submission-materials="true" style="visibility: visible; opacity: 1;" aria-busy="false" data-savescroll="0" aria-hidden="true"><div jsname="a9kxte" class="T4LgNb "><div jsname="qJTHM" class="kFwPee"><div class="xgkURe mhCMAe"></div><div class="xgkURe ECPFEb"></div><div jsaction="rcuQ6b:rcuQ6b" jscontroller="FRimSc"></div><div jscontroller="UqV0cb" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b"><div jscontroller="cs6ocd" jsaction="rcuQ6b:npT2md;FttMgb:Qp7hp;qFdNBb:Pb2hxc;Cvbxce:N6n54b;mlnRJb:p5Uonb" style="display: none;" data-wait-for="QlRoyd"></div><div class="fJ1Vac"><div class="P47N4e vUBwW m1PbN bFjUmb-Wvd9Cc pOf0gc"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M7 15h7v2H7zm0-4h10v2H7zm0-4h10v2H7z"></path><path d="M19 3h-4.18C14.4 1.84 13.3 1 12 1c-1.3 0-2.4.84-2.82 2H5c-.14 0-.27.01-.4.04a2.008 2.008 0 0 0-1.44 1.19c-.1.23-.16.49-.16.77v14c0 .27.06.54.16.78s.25.45.43.64c.27.27.62.47 1.01.55.13.02.26.03.4.03h14c1.1 0 2-.9 2-2V5c0-1.1-.9-2-2-2zm-7-.25c.41 0 .75.34.75.75s-.34.75-.75.75-.75-.34-.75-.75.34-.75.75-.75zM19 19H5V5h14v14z"></path></svg></div><div class="EE538" role="main"><div jscontroller="QlRoyd" jsmodel="I8BbUd;UvJ3Mb;uJydvc;xeYtDf;" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;wJx4ze:rcuQ6b"><div class="nl5VRd ypv4re"><div class="N5dSp"><h1 class="fOvfyc B7SYid VnOHwf-Tvm9db"><span style="white-space: pre-wrap;">LAB03</span></h1><div class="Nmpzvc"></div><div jscontroller="bkcTxe" jsmodel="I8BbUd;PTCFbe" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;wJx4ze:rcuQ6b;aWRkAb:yG0upc" data-hide-copy-link="false" data-hide-delete="false" data-stream-item-id="543303401379" class="I0naMd"><div jsshadow="" role="button" class="U26fgb JRtysb WzwrXb I12f0b K2mXPb wwnMtb oxacD" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" jsname="LgbsSe" tabindex="0" aria-haspopup="true" aria-expanded="false" data-dynamic="true" data-alignright="true" aria-label="Opções de atividades"><div class="NWlf3e MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="MhXXcc oJeWuf"><span class="Lw7GHd snByac"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 8c1.1 0 2-.9 2-2s-.9-2-2-2-2 .9-2 2 .9 2 2 2zm0 2c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2zm0 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2z"></path></svg></span></span></div></div></div><div class="rec5Nb cSyPgb QRiHXd"><div class="YVvGBb">Ricardo Pannain</div><div class="DwLQSc" aria-hidden="true">•</div><div class="YVvGBb">8 de mar.&nbsp;Editado às 21 de mar.</div></div><div class="W4hhKd"><div class="CzuI5c asQXV QRiHXd"><div class="YVvGBb"><div jsaction="rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b" jscontroller="teDhve">100 pontos</div></div></div><div class="asQXV hnID5d"></div></div><div class="Wa3mee nQaZq"><div jscontroller="IGT0cf" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;JIbuQc:Yh7j1c(PlbUX)" jsmodel="xvu37b" data-type="2" data-visibility="2" guidedhelpid="commentsdialogGH" class=" LhPqk" data-with-icon="true" data-show-add-comments-link="true"><div role="button" class="uArJ5e cd29Sd UQuaGc kCyAyd oxacD" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;" jsshadow="" jsname="PlbUX" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue cd29Sd"><span class="E6FpNe Ce1Y1c"><svg width="24" height="24" viewBox="0 0 24 24" focusable="false" class=" NMm5M hhikbc"><path d="M21.99 4c0-1.1-.89-2-1.99-2H4c-1.1 0-2 .9-2 2v12c0 1.1.9 2 2 2h14l4 4-.01-18zM4 16V4h16v12H4z"></path><path d="M6 12h12v2H6zm0-3h12v2H6zm0-3h12v2H6z"></path></svg></span><span class="NPEfkd RveJvd snByac"> 2 comentários da turma</span></span></div></div></div></div></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;wuANJc:.CLIENT;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel="PTCFbe hGbFme BrMJ0e" data-is-edit-mode="false" data-filter="0" data-material-parent-id="PTCFbe" data-include-stream-item-materials="true"><div jsname="UYewLd" class="AgzMgb hjqfGd" style=""><div class="MlZb9c xLFtvb " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;IKzbTb:Yo3LPb;wuANJc:.CLIENT" jsname="C2Qrw" data-parent-id="PTCFbe" data-mode="1" data-copies-only="false" data-show-originality-analyses="false" data-forms-only="false" data-read-only="false"><div data-dom-id="18i9CsuLStFUe1Po7bEnQDuZ-XjezSzRC-0-3-2-PDF-lab03_v2023.1.pdf-$2-false-false-false-false-$-$-https://drive.google.com/file/d/18i9CsuLStFUe1Po7bEnQDuZ-XjezSzRC/view?usp=drive_web&amp;authuser=0" class="t2wIBc"><div class="r0VQac QRiHXd Aopndd " jsname="HzV7m" jsaction="JIbuQc:Rsbfue(Rsbfue);"><a class="vwNuXe JkIgWb QRiHXd MymH0d maXJsd" target="_blank" aria-label="Anexo: PDF: lab03_v2023.1.pdf" jsaction="LWntbc" href="https://drive.google.com/file/d/18i9CsuLStFUe1Po7bEnQDuZ-XjezSzRC/view?usp=drive_web&amp;authuser=0" title="lab03_v2023.1.pdf" data-focus-id="hSRGPd-auswjd-18i9CsuLStFUe1Po7bEnQDuZ-XjezSzRC-https://drive.google.com/file/d/18i9CsuLStFUe1Po7bEnQDuZ-XjezSzRC/view?usp=drive_web&amp;authuser=0" data-attachment-id="18i9CsuLStFUe1Po7bEnQDuZ-XjezSzRC"><div class="bxp7vf bHOAdb Niache"><img jsname="q4uQmd" jsaction="error:dyBsCf" class=" " src="dec2_to_4_files/lab03_v2023.1.pdf.png" aria-hidden="true" role="presentation" data-mime-type="application/pdf" data-iml="579593"></div><div class="MM30Lb"><div class="A6dC2c QDKOcc VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">lab03_v2023.1.pdf</div><div class="cSyPgb WInaFd QRiHXd"><div class="QRiHXd"><div class="kRYv9b YVvGBb">PDF</div></div></div></div></a><div class="ZgfM9 QRiHXd"></div></div></div><div data-dom-id="1zQi_4uZTu5Wns9qt6FGTOfJEF6uQsY81-1-3-2-Arquivo compactado-lab03_material_v2023.1.rar-$2-false-false-false-false-$-$-https://drive.google.com/file/d/1zQi_4uZTu5Wns9qt6FGTOfJEF6uQsY81/view?usp=drive_web&amp;authuser=0" class="t2wIBc"><div class="r0VQac QRiHXd Aopndd " jsname="HzV7m" jsaction="JIbuQc:Rsbfue(Rsbfue);"><a class="vwNuXe JkIgWb QRiHXd MymH0d maXJsd" target="_blank" aria-label="Anexo: Arquivo compactado: lab03_material_v2023.1.rar" jsaction="LWntbc" href="https://drive.google.com/file/d/1zQi_4uZTu5Wns9qt6FGTOfJEF6uQsY81/view?usp=drive_web&amp;authuser=0" title="lab03_material_v2023.1.rar" data-focus-id="hSRGPd-auswjd-1zQi_4uZTu5Wns9qt6FGTOfJEF6uQsY81-https://drive.google.com/file/d/1zQi_4uZTu5Wns9qt6FGTOfJEF6uQsY81/view?usp=drive_web&amp;authuser=0" data-attachment-id="1zQi_4uZTu5Wns9qt6FGTOfJEF6uQsY81"><div class="bxp7vf bHOAdb Niache"><img jsname="q4uQmd" jsaction="error:dyBsCf" class=" " src="dec2_to_4_files/logo_drive_2020q4_color_1x_web_48dp.png" aria-hidden="true" role="presentation" data-mime-type="application/x-rar" data-iml="579316"></div><div class="MM30Lb"><div class="A6dC2c QDKOcc VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">lab03_material_v2023.1.rar</div><div class="cSyPgb WInaFd QRiHXd"><div class="QRiHXd"><div class="kRYv9b YVvGBb">Arquivo compactado</div></div></div></div></a><div class="ZgfM9 QRiHXd"></div></div></div><div data-dom-id="1pkcg2xgbtspjpsNRyqr8Vkam6RAjA9Wx-2-3-2-Arquivo compactado-lab03_material_v2023.1.zip-$2-false-false-false-false-$-$-https://drive.google.com/file/d/1pkcg2xgbtspjpsNRyqr8Vkam6RAjA9Wx/view?usp=drive_web&amp;authuser=0" class="t2wIBc"><div class="r0VQac QRiHXd Aopndd " jsname="HzV7m" jsaction="JIbuQc:Rsbfue(Rsbfue);"><a class="vwNuXe JkIgWb QRiHXd MymH0d maXJsd" target="_blank" aria-label="Anexo: Arquivo compactado: lab03_material_v2023.1.zip" jsaction="LWntbc" href="https://drive.google.com/file/d/1pkcg2xgbtspjpsNRyqr8Vkam6RAjA9Wx/view?usp=drive_web&amp;authuser=0" title="lab03_material_v2023.1.zip" data-focus-id="hSRGPd-auswjd-1pkcg2xgbtspjpsNRyqr8Vkam6RAjA9Wx-https://drive.google.com/file/d/1pkcg2xgbtspjpsNRyqr8Vkam6RAjA9Wx/view?usp=drive_web&amp;authuser=0" data-attachment-id="1pkcg2xgbtspjpsNRyqr8Vkam6RAjA9Wx"><div class="bxp7vf bHOAdb Niache"><img jsname="q4uQmd" jsaction="error:dyBsCf" class=" " src="dec2_to_4_files/logo_drive_2020q4_color_1x_web_48dp.png" aria-hidden="true" role="presentation" data-mime-type="application/x-zip-compressed" data-iml="579316"></div><div class="MM30Lb"><div class="A6dC2c QDKOcc VBEdtc-Wvd9Cc zZN2Lb-Wvd9Cc">lab03_material_v2023.1.zip</div><div class="cSyPgb WInaFd QRiHXd"><div class="QRiHXd"><div class="kRYv9b YVvGBb">Arquivo compactado</div></div></div></div></a><div class="ZgfM9 QRiHXd"></div></div></div></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="MlZb9c xLFtvb " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="1" data-material-parent-id="PTCFbe"></div></div></div><div jsname="QkPyvd" class="" style="display: none;"></div></div><div jsmodel="WuwnAd;jmgIWd;" jscontroller="F37rhb" jsaction="rcuQ6b:rcuQ6b;LSbPUe:rcuQ6b;voP7ud:rcuQ6b" data-course-id="541235264749" class="Z3wmOd lLBkgb" data-allow-rubric-scoring="false"></div><div class="smtc7c"><div class="GWZ7yf AJFihd LBlAUc YkTkoe"><div class="Dy8Cxc QRiHXd"><span class="z3vRcc">Seus trabalhos<div jscontroller="FQo2Xb" jsaction="rcuQ6b:hDYvKe;voP7ud:hDYvKe;qFdNBb:Pb2hxc"></div></span><span class="asQXV"><span jsaction="rcuQ6b:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;uwjiC:rcuQ6b" jscontroller="o5ZA8b" class="UhYXkc KI1A1e ZnNi8e" data-submission-id="2" data-render-simple-labels="true"><span class="u7S8tc YVvGBb"><span class="vzcr8">Atribuído</span></span><span class="E70Hue neggzd" aria-hidden="true">Estigfend</span></span></span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel=" hGbFme BrMJ0e" data-is-edit-mode="false" data-filter="1" data-material-parent-id="2"><div jsname="UYewLd" class="AgzMgb " style="display: none;"><div jscontroller="KqB22e" jsmodel="I8BbUd;PTCFbe;" data-include-stream-item-materials="true" jsaction="rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;mbUMkc:rcuQ6b;IKzbTb:Yo3LPb;wJx4ze:rcuQ6b" jsname="C2Qrw" class="CG2qQ P2wHlc" style="display: none;"></div><div class="JY4wBc MlZb9c " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;IKzbTb:Yo3LPb" jsname="C2Qrw" data-parent-id="2" data-mode="6" data-copies-only="false" data-show-originality-analyses="true" data-forms-only="false" data-read-only="false"></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="JY4wBc MlZb9c " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="6" data-material-parent-id="2"></div></div></div><div jsname="QkPyvd" class="Jp15We tLDEHd B2pRjc" style="">Nenhum trabalho anexado</div><div class="IPGLSb"><div class="QRiHXd J2Cevf" guidedhelpid="submissionManager"><div jsaction="rcuQ6b:rcuQ6b;ln5gI:rcuQ6b;RwVyRc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:rcuQ6b;LEpEAf:qRU3cb" jscontroller="PykWJd" jsmodel="AKq4rd" data-user-id="30751363934" data-attach-actions-control-type="3" data-parent-id="2" class="TDK0Zb CG2qQ cYYbdd"><div jsshadow="" role="button" class="U26fgb REtOWc cd29Sd p0oLxb BEAGS" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" aria-disabled="false" tabindex="0" aria-haspopup="true" aria-expanded="false" guidedhelpid="addOrCreateMaterial" data-menu-type="3" id="ow1044" __is_owner="true"><div class="bnqxkd MbhUzd" jsname="ksKsZd"></div><div class="GJYBjd CeoRYc" aria-hidden="true"></div><span jsslot="" class="GcVcmc Fxmcue cd29Sd"><span class="lRRqZc Ce1Y1c"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="a7AG0 NMm5M"><path d="M20 13h-7v7h-2v-7H4v-2h7V4h2v7h7v2z"></path></svg></span><span class="RdyDwe snByac">Adicionar ou criar</span></span><div jsname="xl07Ob" style="display: none;" aria-hidden="true"><div role="menu" tabindex="0" class="JPdR6b e5Emjc hVNH5c" jscontroller="uY3Nvd" jsaction="IpSVtb:TvD9Pc;fEN2Ze:xzS4ub;frq95c:LNeFm;cFpp9e:J9oOtd; click:H8nU8b; mouseup:H8nU8b; keydown:I481le; keypress:Kr2w4b; blur:O22p3e; focus:H8nU8b"><div class="XvhY1d" jsaction="mousedown:p8EH2c; touchstart:p8EH2c"><div class="JAPqpe K0NPx"><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Google Drive" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg enable-background="new 0 0 24 24" focusable="false" height="24" viewBox="0 0 24 24" width="24" class="zAg7wc xSP5ic NMm5M"><rect fill="none" height="24" width="24"></rect><path d="M14.35,2.5h-4.7c-0.71,0-1.37,0.38-1.73,0.99L1.58,14.4c-0.36,0.62-0.36,1.38-0.01,2l2.35,4.09c0.36,0.62,1.02,1,1.73,1 h12.68c0.72,0,1.38-0.38,1.73-1l2.35-4.09c0.36-0.62,0.35-1.38-0.01-2L16.08,3.49C15.72,2.88,15.06,2.5,14.35,2.5z M18.34,19.5H5.66 l-2.35-4.09L9.65,4.5h4.7l6.34,10.91L18.34,19.5z M12.9,7.75h-1.8l-4.58,7.98L7.25,17h9.5l0.73-1.27L12.9,7.75z M9.25,15L12,10.2 l2.75,4.8H9.25z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:pau0Hb" data-type="2"><div class="jO7h3c">Google Drive</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Link" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="zAg7wc xSP5ic NMm5M"><path d="M3.9 12c0-1.71 1.39-3.1 3.1-3.1h4V7H7c-2.76 0-5 2.24-5 5s2.24 5 5 5h4v-1.9H7c-1.71 0-3.1-1.39-3.1-3.1zM8 13h8v-2H8v2zm9-6h-4v1.9h4c1.71 0 3.1 1.39 3.1 3.1s-1.39 3.1-3.1 3.1h-4V17h4c2.76 0 5-2.24 5-5s-2.24-5-5-5z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:VORrnc"><div class="jO7h3c">Link</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Arquivo" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="zAg7wc xSP5ic NMm5M"><path d="M15.5 6v10.5c0 2.21-1.79 4-4 4s-4-1.79-4-4V6a2.5 2.5 0 0 1 5 0v9.5c0 .55-.45 1-1 1s-1-.45-1-1V6H9v9.5a2.5 2.5 0 0 0 5 0V6c0-2.21-1.79-4-4-4S6 3.79 6 6v10.5c0 3.04 2.46 5.5 5.5 5.5s5.5-2.46 5.5-5.5V6h-1.5z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:pau0Hb" data-type="1"><div class="jO7h3c">Arquivo</div></div></span><div role="separator" aria-hidden="true" class="kCtYwe"></div><h3 class="mMfeif ubvFYc dDKhVc-Wvd9Cc">Criar novo</h3><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Documentos" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="XxyAsb"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="1"><div class="jO7h3c">Documentos</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Apresentações" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="qurv4d"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="3"><div class="jO7h3c">Apresentações</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Planilhas" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="teCq2b"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="2"><div class="jO7h3c">Planilhas</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Desenhos" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="O1YELb"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="6"><div class="jO7h3c">Desenhos</div></div></span></div></div></div></div></div></div></div><div jscontroller="Glz2Ld" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;JIbuQc:f2nbFb" data-submission-id="2"></div><div jscontroller="krEUN" jsaction="JIbuQc:sFeBqf(sFeBqf),ReqGfd(ReqGfd);rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;nK3Vsc:rcuQ6b;ZQcBrc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:Yo3LPb;R6l5Vd:UApqrc;LNlWBf:IyXkod" class="CG2qQ kg6ice"><div jsshadow="" role="button" class="uArJ5e TuHiFd UQuaGc Y5sE8d" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="sFeBqf" tabindex="0" guidedhelpid="submissionManager_markAsDone"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Marcar como concluída</span></span></div></div></div></div><div jscontroller="cTy1kf" jsmodel="I8BbUd" jsaction="rcuQ6b:TZH2db;wuANJc:TZH2db;voP7ud:TZH2db;wJx4ze:TZH2db"></div></div><div class="GWZ7yf m8BrFf LBlAUc YkTkoe" guidedhelpid="submissionPrivateComments"><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="3" data-visibility="1" data-submission-id="30751363934" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;wuANJc:lswmYb;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário particular</span></div><div class="amzDAb"><div class="QxGMXc asQXV QRiHXd"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Comentários particulares</span></div><div jsshadow="" role="button" class="uArJ5e UQuaGc kCyAyd l3F1ye Epqnjf xAiME" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="zPiFrf" aria-label="Adicionar comentário para Ricardo Pannain" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Adicionar comentário para Ricardo Pannain</span></span></div></div><div class="Ono85c VvAAB"></div></div></div></div><div class="pOf0gc"><div class="eqqrO"><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="2" data-visibility="2" class="PeGHgb Q8U8uc" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="VYv8If QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">2 comentários para a turma</span></div><div class="amzDAb"><div class="lq45g asQXV QRiHXd"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M15 8c0-1.42-.5-2.73-1.33-3.76.42-.14.86-.24 1.33-.24 2.21 0 4 1.79 4 4s-1.79 4-4 4c-.43 0-.84-.09-1.23-.21-.03-.01-.06-.02-.1-.03A5.98 5.98 0 0 0 15 8zm1.66 5.13C18.03 14.06 19 15.32 19 17v3h4v-3c0-2.18-3.58-3.47-6.34-3.87zM9 6c-1.1 0-2 .9-2 2s.9 2 2 2 2-.9 2-2-.9-2-2-2m0 9c-2.7 0-5.8 1.29-6 2.01V18h12v-1c-.2-.71-3.3-2-6-2M9 4c2.21 0 4 1.79 4 4s-1.79 4-4 4-4-1.79-4-4 1.79-4 4-4zm0 9c2.67 0 8 1.34 8 4v3H1v-3c0-2.66 5.33-4 8-4z"></path></svg></span><span class="asQXV QRiHXd">Comentários da turma</span></div></div><div class="ruTJle VvAAB"><div class="dZVZab"><div jsaction="ym8qYd:u4pxTb" jscontroller="dvgIje" class="wJ76ge TIunU"><div class="QRiHXd pMq3Db"><img class="WqfsMd tkmmwb" aria-hidden="true" alt="" src="dec2_to_4_files/unnamed_003.png" data-iml="578946"><div class="G0rp"><div class="YU7iib"><div><a class="gJItbc asQXV" aria-label="Comentário postado por Natan Rodrigues de Oliveira">Natan Rodrigues de Oliveira</a><span class="T8rTjd">19 de mar.</span></div><div class="thiSD Gh0umc" jsaction="JIbuQc:pODwA(IgWJu)"><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db L8jEMd CMmBPd oxacD qk5dFc kpDQ8" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="IgWJu" aria-label="Responder" tabindex="0" data-tooltip="Responder a este comentário" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M16 10H6.83L9 7.83l1.41-1.41L9 5l-6 6 6 6 1.41-1.41L9 14.17 6.83 12H16c1.65 0 3 1.35 3 3v4h2v-4c0-2.76-2.24-5-5-5z"></path></svg></span></span></div><div class="KYmC8d kpDQ8 CG2qQ"><div jscontroller="RrRSXd" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b" jsmodel="I8BbUd" data-comment-id="543712453681"></div></div></div></div><div class="VSWCL tLDEHd"><span style="white-space: pre-wrap;">Olá, professor. Não encontrei o arquivo lab03_material_v2023.1.zip para pegar a entity definida no texto do lab. Poderia postar aqui o caminho?</span></div></div></div></div></div><div class="dZVZab"><div jsaction="ym8qYd:u4pxTb" jscontroller="dvgIje" class="wJ76ge TIunU"><div class="QRiHXd pMq3Db"><img class="WqfsMd tkmmwb" aria-hidden="true" alt="" src="dec2_to_4_files/unnamed_003.jpg" data-iml="578946"><div class="G0rp"><div class="YU7iib"><div><a class="gJItbc asQXV" aria-label="Comentário postado por Ricardo Pannain">Ricardo Pannain</a><span class="T8rTjd">20 de mar.</span></div><div class="thiSD Gh0umc" jsaction="JIbuQc:pODwA(IgWJu)"><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db L8jEMd CMmBPd oxacD qk5dFc kpDQ8" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="IgWJu" aria-label="Responder" tabindex="0" data-tooltip="Responder a este comentário" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M16 10H6.83L9 7.83l1.41-1.41L9 5l-6 6 6 6 1.41-1.41L9 14.17 6.83 12H16c1.65 0 3 1.35 3 3v4h2v-4c0-2.76-2.24-5-5-5z"></path></svg></span></span></div><div class="KYmC8d kpDQ8 CG2qQ"><div jscontroller="RrRSXd" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b" jsmodel="I8BbUd" data-comment-id="543724853903"></div></div></div></div><div class="VSWCL tLDEHd"><span style="white-space: pre-wrap;">Incluído  lab03_material_v2023.1.zip</span></div></div></div></div></div></div><div jsname="uqYDP" class="XNP4U Gh0umc kpDQ8 CMmBPd"><div jsaction="JIbuQc:npVELd(IgWJu),sFeBqf(M2UYVd);laiNib:H2nWWd;A56Kbc:BU3G2c;EiG6ec:ZQdNEd; keydown:Hq2uPe" jscontroller="bUQrJd"><div class="QRiHXd"><img aria-hidden="true" alt="" class="a5lbif tkmmwb AI7uec" src="dec2_to_4_files/unnamed_007.jpg" data-iml="578946"><div class="a5kY4d cjzpkc-Wvd9Cc QRiHXd yUZA2d"><div class="nxIm7c" jsaction="YqO5N:HRfSZd; keydown:Hq2uPe"><div jsaction="rcuQ6b:rcuQ6b;YFq8g:PqP2y; focus:h06R8" data-role="owner,coteacher,student" data-include-invited="false" jscontroller="r9MpRb" jsname="Ufn6O" jsmodel="LQajt" data-course-id="541235264749"><div class="O98Lj" style=""><div class="bswVrf Lzdwhd-BrZSOd" aria-hidden="true">Adicionar comentário para a turma...</div><div id=":j.t" class="LsqTRb Lzdwhd-AyKMt tgNIJf-Wvd9Cc Yiql6e iTy5c editable" tabindex="0" role="textbox" aria-required="true" aria-multiline="true" aria-label="Adicionar comentário para a turma..." g_editable="true" contenteditable="true"></div></div></div></div><div class="QRiHXd apsLYe "><div jsshadow="" role="button" class="uArJ5e Y5FYJe cjq2Db OZ6W0d T8tcPb RDPZE" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="M2UYVd" aria-label="Postar" aria-disabled="true" tabindex="-1" data-tooltip="Postar" data-tooltip-vertical-offset="-12" data-tooltip-horizontal-offset="0"><div class="PDXc1b MbhUzd" jsname="ksKsZd"></div><span jsslot="" class="XuQwKc"><span class="GmuOkf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M hhikbc"><path d="M2 3v18l20-9L2 3zm2 11l9-2-9-2V6.09L17.13 12 4 17.91V14z"></path></svg></span></span></div></div></div></div></div></div></div></div></div></div><aside class="asCVDb BiaLW" role="complementary"><div class="GWZ7yf AJFihd LBlAUc YkTkoe"><div class="Dy8Cxc QRiHXd"><span class="z3vRcc">Seus trabalhos<div jscontroller="FQo2Xb" jsaction="rcuQ6b:hDYvKe;voP7ud:hDYvKe;qFdNBb:Pb2hxc"></div></span><span class="asQXV"><span jsaction="rcuQ6b:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;uwjiC:rcuQ6b" jscontroller="o5ZA8b" class="UhYXkc KI1A1e ZnNi8e" data-submission-id="2" data-render-simple-labels="true"><span class="u7S8tc YVvGBb"><span class="vzcr8">Atribuído</span></span><span class="E70Hue neggzd" aria-hidden="true">Estigfend</span></span></span></div><div jsaction="rcuQ6b:rcuQ6b;URgETb:rcuQ6b;uwjiC:rcuQ6b;ZQcBrc:rcuQ6b;nK3Vsc:.CLIENT" class="sVNOQ" jscontroller="yP6Lwf" jsmodel=" hGbFme BrMJ0e" data-is-edit-mode="false" data-filter="1" data-material-parent-id="2"><div jsname="UYewLd" class="AgzMgb " style="display: none;"><div jscontroller="KqB22e" jsmodel="I8BbUd;PTCFbe;" data-include-stream-item-materials="true" jsaction="rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;mbUMkc:rcuQ6b;IKzbTb:Yo3LPb;wJx4ze:rcuQ6b" jsname="C2Qrw" class="CG2qQ P2wHlc" style="display: none;"></div><div class="JY4wBc MlZb9c " jscontroller="ze9NU" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;KtPeHe:rcuQ6b;voP7ud:rcuQ6b;wuANJc:rcuQ6b;IKzbTb:Yo3LPb" jsname="C2Qrw" data-parent-id="2" data-mode="6" data-copies-only="false" data-show-originality-analyses="true" data-forms-only="false" data-read-only="false"></div><div jsmodel="xLJwSb" class="F8dn3e"><div class="JY4wBc MlZb9c " jscontroller="Z2vwzc" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;nK3Vsc:hVCa3c;n7J2fb:GDCStd;IKzbTb:M3TAie;YCR7Tc:STeVHc" jsname="C2Qrw" data-mode="6" data-material-parent-id="2"></div></div></div><div jsname="QkPyvd" class="Jp15We tLDEHd B2pRjc" style="">Nenhum trabalho anexado</div><div class="IPGLSb"><div class="QRiHXd J2Cevf" guidedhelpid="submissionManager"><div jsaction="rcuQ6b:rcuQ6b;ln5gI:rcuQ6b;RwVyRc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:rcuQ6b;LEpEAf:qRU3cb" jscontroller="PykWJd" jsmodel="AKq4rd" data-user-id="30751363934" data-attach-actions-control-type="3" data-parent-id="2" class="TDK0Zb CG2qQ cYYbdd"><div jsshadow="" role="button" class="U26fgb REtOWc cd29Sd p0oLxb BEAGS" jscontroller="iSvg6e" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue; focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;keydown:I481le" aria-disabled="false" tabindex="0" aria-haspopup="true" aria-expanded="false" guidedhelpid="addOrCreateMaterial" data-menu-type="3"><div class="bnqxkd MbhUzd" jsname="ksKsZd"></div><div class="GJYBjd CeoRYc" aria-hidden="true"></div><span jsslot="" class="GcVcmc Fxmcue cd29Sd"><span class="lRRqZc Ce1Y1c"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="a7AG0 NMm5M"><path d="M20 13h-7v7h-2v-7H4v-2h7V4h2v7h7v2z"></path></svg></span><span class="RdyDwe snByac">Adicionar ou criar</span></span><div jsname="xl07Ob" style="display: none;" aria-hidden="true"><div role="menu" tabindex="0" class="JPdR6b e5Emjc hVNH5c" jscontroller="uY3Nvd" jsaction="IpSVtb:TvD9Pc;fEN2Ze:xzS4ub;frq95c:LNeFm;cFpp9e:J9oOtd; click:H8nU8b; mouseup:H8nU8b; keydown:I481le; keypress:Kr2w4b; blur:O22p3e; focus:H8nU8b"><div class="XvhY1d" jsaction="mousedown:p8EH2c; touchstart:p8EH2c"><div class="JAPqpe K0NPx"><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Google Drive" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg enable-background="new 0 0 24 24" focusable="false" height="24" viewBox="0 0 24 24" width="24" class="zAg7wc xSP5ic NMm5M"><rect fill="none" height="24" width="24"></rect><path d="M14.35,2.5h-4.7c-0.71,0-1.37,0.38-1.73,0.99L1.58,14.4c-0.36,0.62-0.36,1.38-0.01,2l2.35,4.09c0.36,0.62,1.02,1,1.73,1 h12.68c0.72,0,1.38-0.38,1.73-1l2.35-4.09c0.36-0.62,0.35-1.38-0.01-2L16.08,3.49C15.72,2.88,15.06,2.5,14.35,2.5z M18.34,19.5H5.66 l-2.35-4.09L9.65,4.5h4.7l6.34,10.91L18.34,19.5z M12.9,7.75h-1.8l-4.58,7.98L7.25,17h9.5l0.73-1.27L12.9,7.75z M9.25,15L12,10.2 l2.75,4.8H9.25z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:pau0Hb" data-type="2"><div class="jO7h3c">Google Drive</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Link" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="zAg7wc xSP5ic NMm5M"><path d="M3.9 12c0-1.71 1.39-3.1 3.1-3.1h4V7H7c-2.76 0-5 2.24-5 5s2.24 5 5 5h4v-1.9H7c-1.71 0-3.1-1.39-3.1-3.1zM8 13h8v-2H8v2zm9-6h-4v1.9h4c1.71 0 3.1 1.39 3.1 3.1s-1.39 3.1-3.1 3.1h-4V17h4c2.76 0 5-2.24 5-5s-2.24-5-5-5z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:VORrnc"><div class="jO7h3c">Link</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Arquivo" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class="zAg7wc xSP5ic NMm5M"><path d="M15.5 6v10.5c0 2.21-1.79 4-4 4s-4-1.79-4-4V6a2.5 2.5 0 0 1 5 0v9.5c0 .55-.45 1-1 1s-1-.45-1-1V6H9v9.5a2.5 2.5 0 0 0 5 0V6c0-2.21-1.79-4-4-4S6 3.79 6 6v10.5c0 3.04 2.46 5.5 5.5 5.5s5.5-2.46 5.5-5.5V6h-1.5z"></path></svg></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:pau0Hb" data-type="1"><div class="jO7h3c">Arquivo</div></div></span><div role="separator" aria-hidden="true" class="kCtYwe"></div><h3 class="mMfeif ubvFYc dDKhVc-Wvd9Cc">Criar novo</h3><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Documentos" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="XxyAsb"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="1"><div class="jO7h3c">Documentos</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Apresentações" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="qurv4d"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="3"><div class="jO7h3c">Apresentações</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Planilhas" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="teCq2b"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="2"><div class="jO7h3c">Planilhas</div></div></span><span jsslot="" jsname="j7LFlb" tabindex="-1" class="z80M1 FeRvI rkHJle" jsaction="click:o6ZaF(preventDefault=true); mousedown:lAhnzb; mouseup:Osgxgf; mouseenter:SKyDAe; mouseleave:xq3APb;touchstart:jJiBRc; touchmove:kZeBdd; touchend:VfAz8(preventMouseEvents=true)" aria-label="Desenhos" role="menuitem"><div class="aBBjbd MbhUzd" jsname="ksKsZd"></div><div class="PCdOIb Ce1Y1c" aria-hidden="true"><div class="O1YELb"></div></div><div class="uyYuVb oJeWuf" jsaction="JIbuQc:v9F4Yd" data-type="6"><div class="jO7h3c">Desenhos</div></div></span></div></div></div></div></div></div></div><div jscontroller="Glz2Ld" jsaction="rcuQ6b:rcuQ6b;uwjiC:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;JIbuQc:f2nbFb" data-submission-id="2"></div><div jscontroller="krEUN" jsaction="JIbuQc:sFeBqf(sFeBqf),ReqGfd(ReqGfd);rcuQ6b:rcuQ6b;wuANJc:rcuQ6b;voP7ud:rcuQ6b;qxfl9d:rcuQ6b;nK3Vsc:rcuQ6b;ZQcBrc:rcuQ6b;uwjiC:rcuQ6b;IKzbTb:Yo3LPb;R6l5Vd:UApqrc;LNlWBf:IyXkod" class="CG2qQ kg6ice"><div jsshadow="" role="button" class="uArJ5e TuHiFd UQuaGc Y5sE8d" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="sFeBqf" tabindex="0" guidedhelpid="submissionManager_markAsDone"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Marcar como concluída</span></span></div></div></div></div><div jscontroller="cTy1kf" jsmodel="I8BbUd" jsaction="rcuQ6b:TZH2db;wuANJc:TZH2db;voP7ud:TZH2db;wJx4ze:TZH2db"></div></div><div class="GWZ7yf m8BrFf LBlAUc YkTkoe" guidedhelpid="submissionPrivateComments"><div jscontroller="XGZuGb" jsmodel="xvu37b;I8BbUd;uJydvc;BCjFBc;" data-type="3" data-visibility="1" data-submission-id="30751363934" class="PeGHgb" jsaction="rcuQ6b:rcuQ6b;Ts0WYd:rcuQ6b;wJx4ze:rcuQ6b;uwjiC:rcuQ6b;wuANJc:lswmYb;JIbuQc:NZUzf(zPiFrf)"><div jsname="tJHJj" jsaction="JIbuQc:jkaCtf" class="WuChGe QRiHXd aHTZpf"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Nenhum comentário particular</span></div><div class="amzDAb"><div class="QxGMXc asQXV QRiHXd"><span class="xSP5ic ho6Zoe bxp7vf"><svg focusable="false" width="24" height="24" viewBox="0 0 24 24" class=" NMm5M"><path d="M12 6c1.1 0 2 .9 2 2s-.9 2-2 2-2-.9-2-2 .9-2 2-2m0 9c2.7 0 5.8 1.29 6 2v1H6v-.99c.2-.72 3.3-2.01 6-2.01m0-11C9.79 4 8 5.79 8 8s1.79 4 4 4 4-1.79 4-4-1.79-4-4-4zm0 9c-2.67 0-8 1.34-8 4v3h16v-3c0-2.66-5.33-4-8-4z"></path></svg></span><span class="asQXV QRiHXd">Comentários particulares</span></div><div jsshadow="" role="button" class="uArJ5e UQuaGc kCyAyd l3F1ye Epqnjf xAiME" jscontroller="VXdfxd" jsaction="click:cOuCgd; mousedown:UX7yZ; mouseup:lbsD7e; mouseenter:tfO1Yc; mouseleave:JywGue;touchstart:p6p2H; touchmove:FwuNnf; touchend:yfqBxc(preventMouseEvents=true|preventDefault=true); touchcancel:JMtRjd;focus:AHmuwe; blur:O22p3e; contextmenu:mg9Pef" jsname="zPiFrf" aria-label="Adicionar comentário para Ricardo Pannain" tabindex="0"><div class="Fvio9d MbhUzd" jsname="ksKsZd"></div><div class="e19J0b CeoRYc"></div><span jsslot="" class="l4V7wb Fxmcue"><span class="NPEfkd RveJvd snByac">Adicionar comentário para Ricardo Pannain</span></span></div></div><div class="Ono85c VvAAB"></div></div></div></aside></div></div><div jscontroller="rFwfKe" jsaction="qFdNBb:Pb2hxc;pN3Oaf:n3lXYe;uwjiC:T0iadd;wuANJc:T0iadd;voP7ud:T0iadd"></div><div jscontroller="BbOAsf" jsmodel="PTCFbe;" jsaction="qFdNBb:Pb2hxc;Cvbxce:ysXIce;pN3Oaf:n3lXYe;wuANJc:hDYvKe,T0iadd;ywGDo:hDYvKe;rcuQ6b:npT2md" data-include-stream-item-materials="true" data-with-stream-item-materials=""></div><div jsaction="Cvbxce:ysXIce;qFdNBb:Pb2hxc;uwjiC:xtpvtf;rcuQ6b:npT2md" jscontroller="cpx3"></div><div jsaction="rcuQ6b:OuAj6c;uwjiC:OuAj6c" jscontroller="ZlX84d" id="ow994" __is_owner="true"></div></div></div><c-data id="c20"></c-data><view-header style="display: none;"><title>Detalhes da atividade</title></view-header></c-wiz><div class="ndfHFb-c4YZDc ndfHFb-c4YZDc-AHmuwe-Hr88gd-OWB6Me dif24c XV0XSd LgGVmb bvmRsc ndfHFb-c4YZDc-vyDMJf-aZ2wEe ndfHFb-c4YZDc-i5oIFb ndfHFb-c4YZDc-TSZdd" aria-label="Mostrando leitor." role="dialog" tabindex="0"><div class="ndfHFb-c4YZDc-bnBfGc ndfHFb-c4YZDc-zTETae" tabindex="0" aria-label="Exibindo lab03_v2023.1.pdf…"></div><div class="ndfHFb-c4YZDc-JNEHMb"></div><div class="ndfHFb-c4YZDc-K9a4Re" style="bottom: 0px; top: 0px;"><div class="ndfHFb-c4YZDc-E7ORLb-LgbsSe ndfHFb-c4YZDc-LgbsSe-OWB6Me ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; left: 12px; opacity: 1;" aria-disabled="true" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="r,c" data-tooltip-offset="-6"><div class="ndfHFb-c4YZDc-DH6Rkf-AHe6Kc"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-tJiF1e-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; right: 12px; opacity: 1;" aria-disabled="false" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="l,c" data-tooltip-offset="-6" tabindex="0" aria-label="Próximo" data-tooltip="Próximo"><div class="ndfHFb-c4YZDc-DH6Rkf-AHe6Kc"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-q77wGc" style="opacity: 1;"><div class="ndfHFb-c4YZDc-DARUcf-NnAfwf-i5oIFb" style="" aria-label="Página 4 de 6"><div class="ndfHFb-c4YZDc-DARUcf-NnAfwf-tJHJj">Página</div><div class="ndfHFb-c4YZDc-DARUcf-NnAfwf-cQYSPc">4</div><span class="ndfHFb-c4YZDc-DARUcf-NnAfwf-hgDUwe">/</span><div class="ndfHFb-c4YZDc-DARUcf-NnAfwf-j4LONd">6</div></div><div class="ndfHFb-c4YZDc-nJjxad-nK2kYb-i5oIFb" style=""><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-nJjxad-m9bMae-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-LgbsSe-OWB6Me" role="button" style="user-select: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Diminuir o zoom" data-tooltip="Diminuir o zoom" aria-disabled="true"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-nJjxad-hj4D6d-LgbsSe VIpgJd-TzA9Ye-eEGnhe" role="button" style="user-select: none;" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Ajustar à largura" data-tooltip="Ajustar à largura"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-nJjxad-bEDTcc-LgbsSe VIpgJd-TzA9Ye-eEGnhe" role="button" style="user-select: none;" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Aumentar o zoom" data-tooltip="Aumentar o zoom"><div class="ndfHFb-c4YZDc-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-LzGo7c" style="display: none;"></div></div><div class="ndfHFb-c4YZDc-K9a4Re-nKQ6qf ndfHFb-c4YZDc-TvD9Pc-qnnXGd" role="main" style=""><div class="ndfHFb-c4YZDc-EglORb-ge6pde ndfHFb-c4YZDc-K9a4Re-ge6pde-Ne3sFf" role="status" tabindex="-1" aria-label="Carregando" style="display: none;"><div class="ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div><span class="ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" aria-hidden="true">Carregando…</span></div><div style="display:none" id="drive-active-item-info">{"id": "18i9CsuLStFUe1Po7bEnQDuZ-XjezSzRC", "title": "lab03_v2023.1.pdf", "mimeType": "application\/pdf"}</div><div class="ndfHFb-c4YZDc-cYSp0e ndfHFb-c4YZDc-oKVyEf"><textarea class="ndfHFb-c4YZDc-cYSp0e-B7I4Od" aria-hidden="true" tabindex="-1"></textarea><div class="ndfHFb-c4YZDc-cYSp0e-s2gQvd ndfHFb-c4YZDc-s2gQvd ndfHFb-c4YZDc-s2gQvd-sn54Q" tabindex="-1" style="margin-left: 12px;"><div class="ndfHFb-c4YZDc-cYSp0e-Oz6c3e ndfHFb-c4YZDc-cYSp0e-DARUcf-gSKZZ ndfHFb-c4YZDc-neVct-RCfa3e" role="document" tabindex="0" style="margin-top: 56px; margin-bottom: 56px; width: 800px; left: 50px;"><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf" style="padding-bottom: 141.25%;"><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf"><a href="https://forms.gle/pUcMCjhBm7faUMWWA" target="_blank" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-hSRGPd" tabindex="0" role="link" aria-label="https://forms.gle/pUcMCjhBm7faUMWWA" data-saferedirecturl="https://www.google.com/url?q=https://forms.gle/pUcMCjhBm7faUMWWA&amp;sa=D&amp;source=apps-viewer-frontend&amp;ust=1680043280504813&amp;usg=AOvVaw2XePFYUmYiG80d0JDIwE72&amp;hl=pt-BR" rel="noreferrer" style="left: 68.9597%; top: 47.2684%; width: 16.7785%; height: 2.019%;"></a><a href="https://forms.gle/pUcMCjhBm7faUMWWA" target="_blank" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-hSRGPd" tabindex="0" role="link" aria-label="https://forms.gle/pUcMCjhBm7faUMWWA" data-saferedirecturl="https://www.google.com/url?q=https://forms.gle/pUcMCjhBm7faUMWWA&amp;sa=D&amp;source=apps-viewer-frontend&amp;ust=1680043280504901&amp;usg=AOvVaw2atbPEqeQ0POwvfTFTJGRM&amp;hl=pt-BR" rel="noreferrer" style="left: 20.8054%; top: 48.9311%; width: 37.5839%; height: 2.019%;"></a></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf"><h2 class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj" tabindex="0">Página 1 de 6</h2><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 34.396%; top: 9.26366%; width: 31.2081%; height: 1.78147%;">MC613 – Laboratório de Circuitos Lógicos
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 42.1141%; top: 17.8147%; width: 15.4362%; height: 1.78147%;">Laboratório 03
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 20.3088%; width: 11.0738%; height: 1.66271%;">Instruções:
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 23.6342%; width: 68.6242%; height: 1.66271%;">- Quando for demonstrar seu trabalho, tome nota do número da placa
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 25.1781%; width: 64.7651%; height: 1.78147%;">utilizada. O número da placa será utilizado para atribuir a nota ao grupo.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 28.0285%; width: 68.6242%; height: 1.78147%;">- A última página deste documento contém um checklist com todos os
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 29.6912%; width: 33.7248%; height: 1.66271%;">arquivos que fazem parte da entrega.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 32.5416%; width: 68.6242%; height: 1.66271%;">- Os nomes dos arquivos devem ser seguidos, e isso faz parte da
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 34.2043%; width: 9.39597%; height: 1.66271%;">avaliação.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 37.0546%; width: 68.6242%; height: 1.66271%;">- A entrega deverá estar em único arquivo .ZIP, com o nome
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 38.5986%; width: 65.604%; height: 1.78147%;">T_Lab03_RA.zip, T é a turma, e RA é o RA do componente do grupo
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 40.2613%; width: 65.604%; height: 1.66271%;">que fará a entrega. Por exemplo, B_Lab03_123456.zip é a entrega do
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 41.924%; width: 41.7785%; height: 1.66271%;">grupo do aluno com o RA 123456, na turma B.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 44.7744%; width: 56.7114%; height: 1.66271%;">- Não divida ou agrupe em pastas os arquivos dentro do .ZIP.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 47.5059%; width: 68.6242%; height: 1.78147%;">- A entrega deve ser feita pelo Google Forms
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 49.1686%; width: 65.604%; height: 1.78147%;">(https://forms.gle/pUcMCjhBm7faUMWWA). Você deve estar autenticado
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 50.8314%; width: 61.9128%; height: 1.66271%;">com uma conta do Google - pode ser uma conta pessoal ou da DAC.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 53.6817%; width: 53.1879%; height: 1.66271%;">- Apenas um integrante do grupo precisa fazer a entrega.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 56.5321%; width: 68.6242%; height: 1.66271%;">- Preste especial atenção aos nomes das entidades e sinais (entradas e
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 58.076%; width: 63.7584%; height: 1.78147%;">saídas) descritos nos laboratórios. Isso também faz parte da avaliação.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 60.9264%; width: 68.6242%; height: 1.78147%;">- Se mais do que um arquivo for recebido para a mesma entrega, o último
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 62.5891%; width: 62.2483%; height: 1.66271%;">recebido será considerado. Utilize o mesmo RA do aluno entregando.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 65.4394%; width: 68.6242%; height: 1.66271%;">- Faça o download do arquivo lab03_material_v2023.1.zip. Esse arquivo
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 19.9664%; top: 67.1021%; width: 65.7718%; height: 1.66271%;">já contém as descrições de entity necessárias para implementar os
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 20.1342%; top: 68.7649%; width: 33.3893%; height: 1.54394%;">circuitos. Utilize elas, e não as altere.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 91.0926%; width: 15.9396%; height: 1.42518%;">Versão 01/03/2023.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 47.9866%; top: 92.7553%; width: 1.00671%; height: 1.30641%;">1
</p></div><div class="ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q" style="display: none;"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b"></div><img src="blob:https://classroom.google.com/a8840637-8e50-4b69-9ab5-3d053d9a4faa" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c" alt="Página 1 de 6" aria-hidden="true"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf" style="padding-bottom: 141.25%;"><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf"><h2 class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj" tabindex="0">Página 2 de 6</h2><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 34.396%; top: 9.26366%; width: 31.2081%; height: 1.78147%;">MC613 – Laboratório de Circuitos Lógicos
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 38.0873%; top: 15.677%; width: 23.8255%; height: 1.42518%;">Parte I - Crossbar switch
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 19.0024%; width: 71.6443%; height: 1.66271%;">Seja o componente xbar que implementa um crossbar switch
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 20.6651%; width: 71.4765%; height: 1.66271%;">(a inversão só ocorre se o S estiver no no nível lógico alto, ou seja, se S = '1').
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 22.209%; width: 71.6443%; height: 1.78147%;">Projete os circuitos abaixo em VHDL e verifique o funcionamento de todos os
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 23.8717%; width: 21.9799%; height: 1.78147%;">projetos com simulação.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 41.4489%; width: 71.4765%; height: 1.66271%;">I.1. Projete este circuito usando a construção WITH, SELECT e WHEN [sem
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 43.1116%; width: 58.0537%; height: 1.66271%;">usar processo]. Teste por simulação. Salve como xbar_v1.vhd.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 46.3183%; width: 71.4765%; height: 1.78147%;">ENTREGAR: Arquivo xbar_v1.vhd e screenshot da simulação em
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 47.981%; width: 12.7517%; height: 1.78147%;">xbar_v1.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 51.3064%; width: 71.6443%; height: 1.66271%;">I.2. Projete este mesmo circuito usando a construção WHEN ELSE [sem usar
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 52.9691%; width: 53.3557%; height: 1.66271%;">processo]. Teste por simulação. Salve como xbar_v2.vhd.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 56.1758%; width: 71.4765%; height: 1.66271%;">ENTREGAR: Arquivo xbar_v2.vhd e screenshot da simulação em
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 57.8385%; width: 12.7517%; height: 1.66271%;">xbar_v2.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 61.1639%; width: 71.4765%; height: 1.66271%;">I.3. Projete este mesmo circuito em VHDL usando a construção PROCESS.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 62.7078%; width: 42.6175%; height: 1.78147%;">Teste por simulação. Salve como xbar_v3.vhd.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 66.0333%; width: 71.4765%; height: 1.66271%;">ENTREGAR: Arquivo xbar_v3.vhd e screenshot da simulação em
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 67.696%; width: 12.7517%; height: 1.66271%;">xbar_v3.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 71.0214%; width: 71.6443%; height: 1.66271%;">I.4. Instanciando alguma das versões do componente xbar acima, implemente
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 72.5653%; width: 71.6443%; height: 1.78147%;">o circuito abaixo, que implementa um número variável de estágios (utilize os
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 74.228%; width: 58.8926%; height: 1.66271%;">comandos GENERIC e GENERATE). Salve como xbar_gen.vhd.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 84.323%; width: 37.2483%; height: 1.54394%;">VCC = constante 1; GND = constante 0
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 85.867%; width: 33.8926%; height: 1.78147%;">ENTREGAR: Arquivo xbar_gen.vhd.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 91.0926%; width: 15.9396%; height: 1.42518%;">Versão 01/03/2023.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 47.651%; top: 92.7553%; width: 1.51007%; height: 1.30641%;">2
</p></div><div class="ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q" style="display: none;"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b"></div><img src="blob:https://classroom.google.com/dac7f2d6-a9b1-40be-9ce9-eef7bcc5c22e" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c" alt="Página 2 de 6" aria-hidden="true"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf" style="padding-bottom: 141.25%;"><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf"><h2 class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj" tabindex="0">Página 3 de 6</h2><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 34.396%; top: 9.26366%; width: 31.2081%; height: 1.78147%;">MC613 – Laboratório de Circuitos Lógicos
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 15.677%; width: 71.6443%; height: 1.78147%;">I.5. Crie um novo projeto instanciando o componente do item I.4 com 5
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 17.3397%; width: 71.6443%; height: 1.66271%;">estágios. Teste por simulação. Salve como xbar_stage_5.vhd. Programe a
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 19.0024%; width: 71.6443%; height: 1.66271%;">placa para verificar o funcionamento, usando 5 switches – SW(0) até SW(4) - e
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 20.6651%; width: 33.3893%; height: 1.66271%;">um LED, sinal LEDR(0), como saída.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 23.8717%; width: 71.6443%; height: 1.78147%;">ENTREGAR: Arquivo xbar_stage_5.vhd e screenshot da simulação em
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 25.5344%; width: 17.953%; height: 1.66271%;">xbar_stage_5.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 28.8599%; width: 71.6443%; height: 1.66271%;">I.6. Repita I.5 para 8 estágios, ou seja, utilizando SW(0) até SW(7). Salve como
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 30.4038%; width: 17.2819%; height: 1.78147%;">xbar_stage_8.vhd
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 33.7292%; width: 71.6443%; height: 1.66271%;">ENTREGAR: Arquivo xbar_stage_8.vhd e screenshot da simulação em
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 35.3919%; width: 17.953%; height: 1.66271%;">xbar_stage_8.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 91.0926%; width: 15.9396%; height: 1.42518%;">Versão 01/03/2023.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 47.8188%; top: 92.7553%; width: 1.1745%; height: 1.42518%;">3
</p></div><div class="ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q" style="display: none;"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b"></div><img src="blob:https://classroom.google.com/82871ba7-d394-4e05-87ac-3a014295eabb" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c" alt="Página 3 de 6" aria-hidden="true"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf" style="padding-bottom: 141.25%;"><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf"><h2 class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj" tabindex="0">Página 4 de 6</h2><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 34.396%; top: 9.26366%; width: 31.2081%; height: 1.78147%;">MC613 – Laboratório de Circuitos Lógicos
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 39.094%; top: 15.677%; width: 21.8121%; height: 1.66271%;">Parte II - Multiplexador
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 19.0024%; width: 71.6443%; height: 1.78147%;">A figura abaixo mostra um circuito multiplexador 4 para 1 projetado
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 20.6651%; width: 71.4765%; height: 1.78147%;">utilizando-se um decodificador 2 para 4 e portas lógicas. w0..3 são as entradas,
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 22.3278%; width: 71.6443%; height: 1.66271%;">s0..1 os sinais de seleção de entrada, En sinal para ligar e desligar o circuito
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 23.9905%; width: 71.6443%; height: 1.66271%;">(significa que, quando desligado, todas as saídas do decodificador serão iguais
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 25.6532%; width: 71.6443%; height: 1.66271%;">à zero) e f a saída selecionada. Projete os circuitos abaixo em VHDL e
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 27.1972%; width: 56.5436%; height: 1.78147%;">verifique o funcionamento de todos os projetos com simulação.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 24.6644%; top: 68.4086%; width: 52.5168%; height: 1.66271%;">Figura 2: Dec2-4 Figura 3: Lógica extra
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 71.9715%; width: 68.1208%; height: 1.66271%;">II.1. Implemente o decodificador 2 para 4 da Figura 2 [sem usar processo].
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 75.1782%; width: 71.6443%; height: 1.78147%;">ENTREGAR: Implementação em VHDL em dec2_to_4.vhd e screenshot da
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 76.8409%; width: 27.8524%; height: 1.78147%;">simulação em dec2_to_4.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 80.1663%; width: 71.6443%; height: 1.66271%;">II.2. Implemente o circuito dentro da caixa pontilhada na Figura 1, conforme o
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 81.829%; width: 38.5906%; height: 1.66271%;">símbolo da Figura 3 [sem usar processo].
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 85.0356%; width: 71.6443%; height: 1.78147%;">ENTREGAR: Implementação em VHDL em extra_logic.vhd e screenshot da
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 86.6983%; width: 28.6913%; height: 1.66271%;">simulação em extra_logic.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 91.0926%; width: 15.9396%; height: 1.42518%;">Versão 01/03/2023.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 47.651%; top: 92.7553%; width: 1.51007%; height: 1.30641%;">4
</p></div><div class="ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q" style="display: none;"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b"></div><img src="blob:https://classroom.google.com/0e5dff28-5dde-4c9b-89d7-054212cde346" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c" alt="Página 4 de 6" aria-hidden="true"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf" style="padding-bottom: 141.25%;"><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf"><h2 class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj" tabindex="0">Página 5 de 6</h2><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 34.396%; top: 9.26366%; width: 31.2081%; height: 1.78147%;">MC613 – Laboratório de Circuitos Lógicos
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 15.677%; width: 71.3087%; height: 1.78147%;">II.3. Instanciando os circuitos dos itens II.1 e II.2, projete um multiplexador 4:1
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 17.3397%; width: 53.8591%; height: 1.66271%;">como na Figura 1. Tabela de mapeamento do multiplexador:
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.4497%; top: 21.0214%; width: 67.7852%; height: 1.78147%;">Valor binário para a porta sel Saída esperada (porta selecionada)
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 30.3691%; top: 24.3468%; width: 39.094%; height: 1.42518%;">00 d0
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 30.3691%; top: 27.5534%; width: 38.7584%; height: 1.42518%;">01 d1
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 30.3691%; top: 30.8789%; width: 39.094%; height: 1.42518%;">10 d2
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 30.5369%; top: 34.0855%; width: 38.9262%; height: 1.42518%;">11 d3
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 39.4299%; width: 71.6443%; height: 1.78147%;">ENTREGAR: Implementação em VHDL em mux4_to_1.vhd e screenshot da
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 41.0926%; width: 28.5235%; height: 1.66271%;">simulação em mux4_to_1.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 44.4181%; width: 71.4765%; height: 1.66271%;">II.4. Instanciando o circuito do item II.3, implemente um multiplexador 16:1 em
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 45.962%; width: 71.6443%; height: 1.78147%;">VHDL. Lembre-se que o quando o valor da entrada sel for igual a 0000, então a
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 47.6247%; width: 71.6443%; height: 1.78147%;">saída o bit menos significativo da porta data, ou seja data(0); e se sel for 1111,
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 49.2874%; width: 71.6443%; height: 1.66271%;">então a saída será o bit mais significativo, ou seja data(15). Não deve ser
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 50.9501%; width: 71.6443%; height: 1.66271%;">usado processo nem implementado de forma estrutural (utilizando portas
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 52.6128%; width: 7.71812%; height: 1.66271%;">lógicas).
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 55.8195%; width: 71.6443%; height: 1.78147%;">ENTREGAR: Implementação em VHDL em mux16_to_1.vhd e screenshot da
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 57.4822%; width: 29.698%; height: 1.66271%;">simulação em mux16_to_1.png.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 91.0926%; width: 15.9396%; height: 1.42518%;">Versão 01/03/2023.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 47.8188%; top: 92.7553%; width: 1.1745%; height: 1.42518%;">5
</p></div><div class="ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q" style="display: none;"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b"></div><img src="blob:https://classroom.google.com/778f79d8-8f39-4f5b-9549-fdc2ecbf5ba7" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c" alt="Página 5 de 6" aria-hidden="true"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf" style="padding-bottom: 141.25%;"><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-PLDbbf"></div><div class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-bN97Pc-haAclf"><h2 class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-tJHJj" tabindex="0">Página 6 de 6</h2><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 34.396%; top: 9.26366%; width: 31.2081%; height: 1.78147%;">MC613 – Laboratório de Circuitos Lógicos
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 42.6175%; top: 15.7957%; width: 14.5973%; height: 1.54394%;">- ENTREGA -
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 20.4276%; width: 71.6443%; height: 1.66271%;">Entregue um único arquivo comprimido em formato ZIP de nome
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 22.0903%; width: 71.4765%; height: 1.66271%;">T_Lab03_RA.zip, onde RA é o RA do aluno entregando e T é a turma,
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 23.753%; width: 9.0604%; height: 1.42518%;">contendo:
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 26.6033%; width: 47.9866%; height: 1.66271%;">- Arquivos xbar_v1.vhd e xbar_v1.png do item I.1.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 28.9786%; width: 47.9866%; height: 1.78147%;">- Arquivos xbar_v2.vhd e xbar_v2.png do item I.2.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 31.4727%; width: 47.9866%; height: 1.66271%;">- Arquivos xbar_v3.vhd e xbar_v3.png do item I.3.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 33.9667%; width: 34.2282%; height: 1.66271%;">- Arquivo xbar_gen.vhd do item I.4.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 36.342%; width: 58.557%; height: 1.78147%;">- Arquivos xbar_stage_5.vhd e xbar_stage_5.png do item I.5.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 38.8361%; width: 58.557%; height: 1.66271%;">- Arquivos xbar_stage_8.vhd e xbar_stage_8.png do item I.6.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 41.3302%; width: 53.0201%; height: 1.66271%;">- Arquivos dec2_to_4.vhd e dec2_to_4.png do item II.1.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 43.7055%; width: 54.698%; height: 1.78147%;">- Arquivos extra_logic.vhd e extra_logic.png do item II.2.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 46.1995%; width: 54.3624%; height: 1.66271%;">- Arquivos mux4_to_1.vhd e mux4_to_1.png do item II.3.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 17.1141%; top: 48.6936%; width: 56.7114%; height: 1.66271%;">- Arquivos mux16_to_1.vhd e mux16_to_1.png do item II.4.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 14.094%; top: 91.0926%; width: 15.9396%; height: 1.42518%;">Versão 01/03/2023.
</p><p class="ndfHFb-c4YZDc-cYSp0e-DARUcf-Df1ZY-eEGnhe" style="left: 47.8188%; top: 92.7553%; width: 1.34228%; height: 1.42518%;">6
</p></div><div class="ndfHFb-c4YZDc-cYSp0e-wxLEad-sn54Q" style="display: none;"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-gvZm2b"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-vWsuo-fmcmS-G0jgYd"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-IDNFyf ndfHFb-c4YZDc-cYSp0e-oYxtQd-gvZm2b"></div><img src="blob:https://classroom.google.com/69dbf5e6-da0b-47ed-b68d-3fa5de9b5b7c" class="ndfHFb-c4YZDc-cYSp0e-DARUcf-RJLb9c" alt="Página 6 de 6" aria-hidden="true"></div></div><span class="ndfHFb-c4YZDc-cYSp0e-AznF2e-DTMEae" tabindex="0"></span></div><div class="ndfHFb-c4YZDc-n5VRYe-ma6Yeb" style="display: none;"></div><div class="ndfHFb-c4YZDc-n5VRYe-AeOLfc" style="display: none;"></div><div class="ndfHFb-c4YZDc-n5VRYe-cGMI2b" style="display: none;"></div><div class="ndfHFb-c4YZDc-n5VRYe-hOcTPc" style="display: none;"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe" aria-hidden="true"><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-haAclf"><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf-haAclf"><input class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-YPqjbf V67aGc-YPqjbf-V67aGc" placeholder="Localizar no documento" aria-label="Localizar no documento" tabindex="-1"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf-haAclf"><span class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-NnAfwf"></span></div></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-E7ORLb ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Localizar anterior" data-tooltip="Localizar anterior"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-tJiF1e ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Localizar próximo" data-tooltip="Localizar próximo"></div><div class="ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-TvD9Pc ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-vWsuo-fmcmS-xxlfEe-SKd3Ne VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Fechar barra de pesquisa" data-tooltip="Fechar barra de pesquisa"></div></div></div></div><div class="ndfHFb-c4YZDc-K9a4Re-nKQ6qf ndfHFb-c4YZDc-TvD9Pc-qnnXGd" role="main" style="display: none;"><div class="ndfHFb-c4YZDc-EglORb-ge6pde ndfHFb-c4YZDc-K9a4Re-ge6pde-Ne3sFf" role="status" tabindex="-1" aria-label="Carregando" style=""><div class="ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div><span class="ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" aria-hidden="true">Carregando…</span></div><div style="display:none">{"id": "1zQi_4uZTu5Wns9qt6FGTOfJEF6uQsY81", "title": "lab03_material_v2023.1.rar", "mimeType": "application\/x-rar"}</div><div class="ndfHFb-c4YZDc-oKVyEf ndfHFb-c4YZDc-TvD9Pc-qnnXGd " style="display: none;"><div class="ndfHFb-c4YZDc-oKVyEf-haAclf"><div class="ndfHFb-c4YZDc-s2gQvd ndfHFb-c4YZDc-oKVyEf-s2gQvd"><div class="ndfHFb-c4YZDc-TvD9Pc-qnnXGd"><div class="ndfHFb-c4YZDc-wvGCSb-gkA7Yd"></div></div></div><div class="ndfHFb-c4YZDc-JqEhuc"><div class="ndfHFb-c4YZDc-JqEhuc-tJHJj"><div class="ndfHFb-c4YZDc-JqEhuc-r4nke-tJHJj"><div class="ndfHFb-c4YZDc-JqEhuc-r4nke-oKdM2c"><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-Bz112c"></div><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d" tabindex="-1">Nome</div><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd">Última modificação</div><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe">Tamanho do arquivo</div></div></div><div class="ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6"></div><div class="ndfHFb-c4YZDc-JqEhuc-n5VRYe"></div></div><div class="ndfHFb-c4YZDc-JqEhuc-bN97Pc ndfHFb-c4YZDc-JqEhuc-s2gQvd ndfHFb-c4YZDc-s2gQvd ndfHFb-c4YZDc-s2gQvd-to915 ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae ndfHFb-c4YZDc-S2QgGf-haAclf" aria-label="Lista de conteúdo arquivado " style="user-select: none;" role="listbox" tabindex="0"></div></div></div></div></div><div class="ndfHFb-c4YZDc-K9a4Re-nKQ6qf ndfHFb-c4YZDc-TvD9Pc-qnnXGd" role="main" style="display: none;"><div class="ndfHFb-c4YZDc-EglORb-ge6pde ndfHFb-c4YZDc-K9a4Re-ge6pde-Ne3sFf" role="status" tabindex="-1" aria-label="Carregando" style="display: none;"><div class="ndfHFb-c4YZDc-EglORb-ge6pde-RJLb9c ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div><span class="ndfHFb-c4YZDc-EglORb-ge6pde-fmcmS ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae" aria-hidden="true">Carregando…</span></div><div style="display:none">{"id": "1pkcg2xgbtspjpsNRyqr8Vkam6RAjA9Wx", "title": "lab03_material_v2023.1.zip", "mimeType": "application\/x-zip-compressed"}</div><div class="ndfHFb-c4YZDc-oKVyEf ndfHFb-c4YZDc-TvD9Pc-qnnXGd " style="display: none;"><div class="ndfHFb-c4YZDc-oKVyEf-haAclf"><div class="ndfHFb-c4YZDc-s2gQvd ndfHFb-c4YZDc-oKVyEf-s2gQvd"><div class="ndfHFb-c4YZDc-TvD9Pc-qnnXGd"><div class="ndfHFb-c4YZDc-wvGCSb-gkA7Yd"></div></div></div><div class="ndfHFb-c4YZDc-JqEhuc"><div class="ndfHFb-c4YZDc-JqEhuc-tJHJj"><div class="ndfHFb-c4YZDc-JqEhuc-r4nke-tJHJj"><div class="ndfHFb-c4YZDc-JqEhuc-r4nke-oKdM2c"><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-Bz112c"></div><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-jIkMge-oKdM2c-V1ur5d" tabindex="-1">Nome</div><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-oKdM2c-TzVJe-ihIZgd">Última modificação</div><div class="ndfHFb-c4YZDc-JqEhuc-oKdM2c-dJDgTb ndfHFb-c4YZDc-JqEhuc-oKdM2c-SxQuSe">Tamanho do arquivo</div></div></div><div class="ndfHFb-c4YZDc-JqEhuc-a4fUwd-Bz112c ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6"></div><div class="ndfHFb-c4YZDc-JqEhuc-n5VRYe"></div></div><div class="ndfHFb-c4YZDc-JqEhuc-bN97Pc ndfHFb-c4YZDc-JqEhuc-s2gQvd ndfHFb-c4YZDc-s2gQvd ndfHFb-c4YZDc-s2gQvd-to915 ndfHFb-c4YZDc-AHmuwe-wcotoc-zTETae ndfHFb-c4YZDc-S2QgGf-haAclf" aria-label="Lista de conteúdo arquivado " style="user-select: none;" role="listbox" tabindex="0"></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b" role="toolbar" style="opacity: 1;"><div class="ndfHFb-c4YZDc-Wrql6b-SmKAyb" style="margin-right: 12px; padding-left: 12px;"><div class="ndfHFb-c4YZDc-Wrql6b-hOcTPc" style="left: 12px;"><div class="ndfHFb-c4YZDc-TvD9Pc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Fechar" data-tooltip="Fechar"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div><div class="ndfHFb-c4YZDc-Wrql6b-Bz112c" tabindex="-1" role="img" style="background-image: url(&quot;//ssl.gstatic.com/docs/doclist/images/mediatype/icon_3_pdf_x16.png&quot;); background-position: left top; background-repeat: no-repeat;" aria-label="Ícone de PDF"></div><div class="ndfHFb-c4YZDc-Wrql6b-jfdpUb" tabindex="-1"><div class="ndfHFb-c4YZDc-Wrql6b-V1ur5d" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6">lab03_v2023.1.pdf</div><div class="ndfHFb-c4YZDc-Wrql6b-V1ur5d ndfHFb-c4YZDc-Wrql6b-V1ur5d-hpYHOb">lab03_v2023.1.pdf</div><div class="ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d" style="display: none;"></div><div class="ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d ndfHFb-c4YZDc-Wrql6b-K4efff-V1ur5d-hpYHOb"></div></div><div class="ndfHFb-c4YZDc-Ujd07d-Btuy5e-Bz112c" style="display: none;"></div><div class="ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b"></div></div><div class="ndfHFb-c4YZDc-Wrql6b-DdWCyb-b0t70b" style=""><div class="ndfHFb-c4YZDc-Wrql6b-FNFY6c-J42Xof-qMHh7d" style=""><div class="ndfHFb-c4YZDc-Wrql6b-FNFY6c ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true"><div class="ndfHFb-c4YZDc-FNFY6c-DWWcKd-Bz112c" style="display: none;"></div><div class="ndfHFb-c4YZDc-FNFY6c-V67aGc">Abrir</div></div><div class="ndfHFb-c4YZDc-Wrql6b-PlOyMe ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-Wrql6b-FNFY6c-BP2Omd-qMHh7d" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true"><div class="ndfHFb-c4YZDc-Wrql6b-PlOyMe-bN97Pc">Extrair</div><div class="ndfHFb-c4YZDc-Wrql6b-HDMZaf-Bz112c"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b-qMHh7d ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" aria-expanded="false" aria-haspopup="true" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Abrir com" data-tooltip="Abrir com" aria-hidden="false" tabindex="0"><div class="ndfHFb-c4YZDc-Wrql6b-FNFY6c-hgDUwe"></div><div class="ndfHFb-c4YZDc-Wrql6b-qMHh7d-SmKAyb"><div class="ndfHFb-c4YZDc-Wrql6b-qMHh7d-fmcmS" tabindex="-1">Abrir com</div><div class="ndfHFb-c4YZDc-Wrql6b-xl07Ob-LgbsSe-hFsbo"><div class="ndfHFb-c4YZDc-Bz112c"></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b-zM6fo-GMvhG-b0t70b" style="display: none;"><div class="ndfHFb-c4YZDc-zM6fo-GMvhG-Bz112c ndfHFb-c4YZDc-Bz112c"></div><span class="ndfHFb-c4YZDc-zM6fo-GMvhG-fmcmS" tabindex="0" role="alert"></span></div><div class="ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b"></div></div><div class="ndfHFb-c4YZDc-Wrql6b-AeOLfc-b0t70b"><div class="ndfHFb-c4YZDc-GSQQnc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe" aria-label="Ver em outra janela" style="display: none;"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div><div class="ndfHFb-c4YZDc-Wrql6b-LQLjdd"><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-ndfHFb VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true" aria-label="Adicionar a &quot;Meu Drive&quot;" data-tooltip="Adicionar a &quot;Meu Drive&quot;"><div class="ndfHFb-c4YZDc-Wrql6b-htvI8d-wcotoc-wHEfpf-ndfHFb-Bz112c"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-Wrql6b-C7uZwb-b0t70b"><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-C7uZwb-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-C7uZwb-LgbsSe-SfQLQb-Bz112c" role="button" style="user-select: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-disabled="false" aria-hidden="false" aria-label="Imprimir" data-tooltip="Imprimir" tabindex="0"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c ndfHFb-c4YZDc-PEFSMe-Bz112c"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-C7uZwb-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe ndfHFb-c4YZDc-C7uZwb-LgbsSe-SfQLQb-Bz112c ndfHFb-c4YZDc-LgbsSe-OWB6Me" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-disabled="true" aria-hidden="true" aria-label="Fazer o download" data-tooltip="Fazer o download"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-C7uZwb-LgbsSe-Bz112c ndfHFb-c4YZDc-nupQLb-Bz112c"><div class="ndfHFb-aZ2wEe" dir="ltr"><div class="ndfHFb-vyDMJf-aZ2wEe auswjd"><div class="aZ2wEe-pbTTYe aZ2wEe-v3pZbf"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-oq6NAc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-gS7Ybc"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div><div class="aZ2wEe-pbTTYe aZ2wEe-nllRtd"><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-LK5yu"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-pehrl-TpMipd"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div><div class="aZ2wEe-LkdAo-e9ayKc aZ2wEe-qwU8Me"><div class="aZ2wEe-LkdAo aZ2wEe-hj4D6d"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-z5C9Gb-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe VIpgJd-TzA9Ye-eEGnhe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" aria-expanded="false" aria-haspopup="true" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Mais ações" data-tooltip="Mais ações" aria-hidden="false" tabindex="0"><div class="ndfHFb-c4YZDc-Bz112c"></div></div></div></div></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-b0t70b ndfHFb-c4YZDc-MZArnb-b0t70b-L6cTce" aria-hidden="true"><div class="ndfHFb-c4YZDc-MZArnb-tJHJj"><div class="ndfHFb-c4YZDc-MZArnb-cXCLoc ndfHFb-c4YZDc-MZArnb-cXCLoc-DKlKme ndfHFb-c4YZDc-MZArnb-cXCLoc-ma6Yeb" style="user-select: none;" role="tablist" aria-label="Barra de guias do painel de detalhes. Pressione as teclas de seta esquerda e direita para mudar de guia." aria-activedescendant="dvdt_goog_225443150"><div class="ndfHFb-c4YZDc-MZArnb-AznF2e ndfHFb-c4YZDc-MZArnb-AznF2e-ZmdkE ndfHFb-c4YZDc-MZArnb-AznF2e-gk6SMd" role="tab" style="user-select: none;" aria-selected="true" id="dvdt_goog_225443150" tabindex="0">Detalhes</div><div class="ndfHFb-c4YZDc-MZArnb-AznF2e ndfHFb-c4YZDc-MZArnb-AznF2e-uDEFge" role="tab" style="user-select: none; display: none;" aria-selected="false" id="dvdt_goog_225443151" aria-hidden="true">Comentários</div></div><div class="ndfHFb-c4YZDc-TvD9Pc-LgbsSe ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none;" tabindex="0" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-label="Ocultar detalhes" data-tooltip="Ocultar detalhes"><div class="ndfHFb-c4YZDc-Bz112c ndfHFb-c4YZDc-DH6Rkf-Bz112c"></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-bN97Pc ndfHFb-c4YZDc-s2gQvd"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-nUpftc" role="tabpanel" style="" aria-labelledby="dvdt_goog_225443150"><div role="complementary" aria-label="Informações gerais" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Informações gerais</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-BKwaUc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Tipo</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">PDF</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0" style="display: none;"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Dimensões</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b"></div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Tamanho</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">280 KB</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0" style="display: none;"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Duração</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b"></div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0" style="display: none;"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Local</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b"><div class="ndfHFb-c4YZDc-MZArnb-P86uke-PntVL"></div></div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Modificado</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">09:40 28 de fev.</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Criado</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">07:39 8 de mar.</div></div><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-Tswv1b-V67aGc">Aberto por mim</div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-ibnC6b">19:31 26 de mar.</div></div></div></div></div><div role="complementary" aria-label="Compartilhamento" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Compartilhamento</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-BKwaUc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-V67aGc ndfHFb-c4YZDc-MZArnb-BA389-V67aGc"><div class="ndfHFb-c4YZDc-MZArnb-BA389-YLEF4c"><img class="ndfHFb-c4YZDc-MZArnb-jNm5if-YLEF4c" alt="" src="dec2_to_4_files/unnamed_006.jpg" role="img" data-tooltip="pannain@unicamp.br" aria-label="pannain@unicamp.br" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" data-iml="612735"></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-V1ur5d" data-tooltip="Ricardo Pannain" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" data-tooltip-only-on-overflow="true">Ricardo Pannain</div></div><div class="ndfHFb-c4YZDc-MZArnb-BA389-nNAX0">Proprietário</div></div></div></div></div><div role="complementary" aria-label="Descrição" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Descrição</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true" aria-label="Editar a descrição" data-tooltip="Editar a descrição"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div><div class="ndfHFb-c4YZDc-MZArnb-ij8cu" role="complementary" tabindex="0">Nenhuma descrição</div><textarea class="ndfHFb-c4YZDc-MZArnb-ij8cu-DyVDA ndfHFb-c4YZDc-s2gQvd" role="textbox" aria-multiline="true" style="display: none;"></textarea></div></div></div><div role="complementary" aria-label="Permissão para download" tabindex="-1" style=""><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj"><span class="ndfHFb-c4YZDc-MZArnb-BKwaUc-tJHJj-fmcmS" role="heading">Permissão para download</span><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe-haAclf"><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-hgDUwe"></div></div></div><div class="ndfHFb-c4YZDc-to915-LgbsSe ndfHFb-c4YZDc-MZArnb-DyVDA-LgbsSe ndfHFb-c4YZDc-LgbsSe" role="button" style="user-select: none; display: none;" data-tooltip-unhoverable="true" data-tooltip-delay="500" data-tooltip-class="ndfHFb-c4YZDc-tk3N6e-suEOdc" data-tooltip-align="b,c" data-tooltip-offset="-6" aria-hidden="true"><div class="ndfHFb-c4YZDc-Bz112c"></div></div><div class="ndfHFb-c4YZDc-MZArnb-BKwaUc-bN97Pc"><div class="ndfHFb-c4YZDc-MZArnb-Tswv1b-oKdM2c" tabindex="0"><div class="ndfHFb-c4YZDc-MZArnb-nupQLb-BA389-Ne3sFf" id="dvddp_goog_225443149">Os leitores podem fazer o download</div></div></div></div><div></div><div></div></div><div class="ndfHFb-c4YZDc-MZArnb-RDNXzf-nUpftc" role="tabpanel" style="display: none;" aria-labelledby="dvdt_goog_225443151"></div></div></div></div><span class="ndfHFb-c4YZDc-AznF2e-DTMEae" style="" tabindex="0" aria-hidden="true"></span><iframe id="apiproxy8511870df0af66dda0066b17c8e88495d95cbc950.1262793752" name="apiproxy8511870df0af66dda0066b17c8e88495d95cbc950.1262793752" style="width: 1px; height: 1px; position: absolute; top: -100px; display: none;" src="dec2_to_4_files/proxy.html" tabindex="-1" aria-hidden="true"></iframe><iframe id="apiproxyb3ab305b7f528d2f49fc642f1e845c1f7b7b15220.3572601733" name="apiproxyb3ab305b7f528d2f49fc642f1e845c1f7b7b15220.3572601733" style="width: 1px; height: 1px; position: absolute; top: -100px; display: none;" src="dec2_to_4_files/proxy_002.html" tabindex="-1" aria-hidden="true"></iframe><div class="ndfHFb-c4YZDc-mg9Pef ndfHFb-c4YZDc-mg9Pef-BvBYQ ndfHFb-c4YZDc-i5oIFb" style="user-select: none; display: none;" role="menu" aria-haspopup="true" tabindex="-1" aria-hidden="true"><div class="ndfHFb-c4YZDc-j7LFlb" role="menuitem" style="user-select: none; display: none;" aria-hidden="true" id=":3p"><div class="ndfHFb-c4YZDc-j7LFlb-bN97Pc">Copiar</div></div><div class="ndfHFb-c4YZDc-j7LFlb" role="menuitem" style="user-select: none; display: none;" aria-hidden="true" id=":3q"><div class="ndfHFb-c4YZDc-j7LFlb-bN97Pc">Adicionar um comentário</div></div></div><div id="goog-lr-1097" style="position: absolute; top: -1000px; height: 1px; overflow: hidden;" aria-live="polite" aria-atomic="true">Página 4 de 6</div><div class="ndfHFb-c4YZDc-mg9Pef ndfHFb-c4YZDc-mg9Pef-BvBYQ ndfHFb-c4YZDc-i5oIFb" style="user-select: none; display: none;" role="menu" aria-haspopup="true" tabindex="-1"><div class="ndfHFb-c4YZDc-j7LFlb" role="menuitem" style="user-select: none; display: none;" aria-hidden="true" id=":4u"><div class="ndfHFb-c4YZDc-j7LFlb-bN97Pc">Copiar</div></div><div class="ndfHFb-c4YZDc-j7LFlb" role="menuitem" style="user-select: none; display: none;" aria-hidden="true" id=":4v"><div class="ndfHFb-c4YZDc-j7LFlb-bN97Pc">Adicionar um comentário</div></div></div></body></html>