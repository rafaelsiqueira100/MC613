LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux4_to_1 IS
port(
     	sel[2], en, w : IN STD_LOGIC;
        d0, d1, d2, d3: OUT STD_LOGIC
);
END mux4_to_1;

ARCHITECTURE LogicFunction3 OF mux_4_to_1 IS

BEGIN
     	dec2_to_4
        extra_logic
END;
